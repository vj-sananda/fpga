`define f0_W0_LSB  0
`define f0_W0_MSB  31

`define f1_W1_LSB  0
`define f1_W1_MSB  31

`define f2_W2_LSB  0
`define f2_W2_MSB  31

`define f3_W3_LSB  0
`define f3_W3_MSB  31

`define f4_W4_LSB  0
`define f4_W4_MSB  31

