  assign enable_aim = category_rd[`CATEGORY_aim];
  assign enable_bittorrent = category_rd[`CATEGORY_bittorrent];
  assign enable_cvs = category_rd[`CATEGORY_cvs];
  assign enable_dhcp = category_rd[`CATEGORY_dhcp];
  assign enable_directconnect = category_rd[`CATEGORY_directconnect];
  assign enable_dns = category_rd[`CATEGORY_dns];
  assign enable_fasttrack = category_rd[`CATEGORY_fasttrack];
  assign enable_finger = category_rd[`CATEGORY_finger];
  assign enable_freenet = category_rd[`CATEGORY_freenet];
  assign enable_ftp = category_rd[`CATEGORY_ftp];
  assign enable_gnutella = category_rd[`CATEGORY_gnutella];
  assign enable_gopher = category_rd[`CATEGORY_gopher];
  assign enable_http = category_rd[`CATEGORY_http];
  assign enable_imap = category_rd[`CATEGORY_imap];
  assign enable_irc = category_rd[`CATEGORY_irc];
  assign enable_jabber = category_rd[`CATEGORY_jabber];
  assign enable_msn = category_rd[`CATEGORY_msn];
  assign enable_napster = category_rd[`CATEGORY_napster];
  assign enable_netbios = category_rd[`CATEGORY_netbios];
  assign enable_nntp = category_rd[`CATEGORY_nntp];
  assign enable_pop3 = category_rd[`CATEGORY_pop3];
  assign enable_rlogin = category_rd[`CATEGORY_rlogin];
  assign enable_sip = category_rd[`CATEGORY_sip];
  assign enable_smtp = category_rd[`CATEGORY_smtp];
  assign enable_snmp = category_rd[`CATEGORY_snmp];
  assign enable_socks = category_rd[`CATEGORY_socks];
  assign enable_ssh = category_rd[`CATEGORY_ssh];
  assign enable_ssl = category_rd[`CATEGORY_ssl];
  assign enable_subversion = category_rd[`CATEGORY_subversion];
  assign enable_telnet = category_rd[`CATEGORY_telnet];
  assign enable_tor = category_rd[`CATEGORY_tor];
  assign enable_vnc = category_rd[`CATEGORY_vnc];
  assign enable_worldofwarcraft = category_rd[`CATEGORY_worldofwarcraft];
  assign enable_x11 = category_rd[`CATEGORY_x11];
  assign enable_yahoo = category_rd[`CATEGORY_yahoo];
