`timescale 1ns/1ps

`define ENABLED_REGEX_CATEGORY_napster TRUE

module CATEGORY_napster_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_CATEGORY_napster

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd1;
    1: charMap = 8'd1;
    2: charMap = 8'd2;
    3: charMap = 8'd1;
    4: charMap = 8'd1;
    5: charMap = 8'd1;
    6: charMap = 8'd2;
    7: charMap = 8'd1;
    8: charMap = 8'd1;
    9: charMap = 8'd1;
    10: charMap = 8'd0;
    11: charMap = 8'd1;
    12: charMap = 8'd1;
    13: charMap = 8'd0;
    14: charMap = 8'd1;
    15: charMap = 8'd1;
    16: charMap = 8'd1;
    17: charMap = 8'd1;
    18: charMap = 8'd1;
    19: charMap = 8'd1;
    20: charMap = 8'd1;
    21: charMap = 8'd1;
    22: charMap = 8'd1;
    23: charMap = 8'd1;
    24: charMap = 8'd1;
    25: charMap = 8'd1;
    26: charMap = 8'd1;
    27: charMap = 8'd1;
    28: charMap = 8'd1;
    29: charMap = 8'd1;
    30: charMap = 8'd1;
    31: charMap = 8'd1;
    32: charMap = 8'd4;
    33: charMap = 8'd3;
    34: charMap = 8'd3;
    35: charMap = 8'd3;
    36: charMap = 8'd3;
    37: charMap = 8'd3;
    38: charMap = 8'd3;
    39: charMap = 8'd3;
    40: charMap = 8'd3;
    41: charMap = 8'd3;
    42: charMap = 8'd3;
    43: charMap = 8'd16;
    44: charMap = 8'd3;
    45: charMap = 8'd11;
    46: charMap = 8'd3;
    47: charMap = 8'd3;
    48: charMap = 8'd9;
    49: charMap = 8'd17;
    50: charMap = 8'd13;
    51: charMap = 8'd5;
    52: charMap = 8'd5;
    53: charMap = 8'd5;
    54: charMap = 8'd5;
    55: charMap = 8'd5;
    56: charMap = 8'd5;
    57: charMap = 8'd10;
    58: charMap = 8'd3;
    59: charMap = 8'd3;
    60: charMap = 8'd3;
    61: charMap = 8'd3;
    62: charMap = 8'd3;
    63: charMap = 8'd3;
    64: charMap = 8'd3;
    65: charMap = 8'd3;
    66: charMap = 8'd3;
    67: charMap = 8'd3;
    68: charMap = 8'd3;
    69: charMap = 8'd3;
    70: charMap = 8'd3;
    71: charMap = 8'd3;
    72: charMap = 8'd3;
    73: charMap = 8'd3;
    74: charMap = 8'd3;
    75: charMap = 8'd3;
    76: charMap = 8'd3;
    77: charMap = 8'd3;
    78: charMap = 8'd3;
    79: charMap = 8'd3;
    80: charMap = 8'd3;
    81: charMap = 8'd3;
    82: charMap = 8'd3;
    83: charMap = 8'd3;
    84: charMap = 8'd3;
    85: charMap = 8'd3;
    86: charMap = 8'd3;
    87: charMap = 8'd3;
    88: charMap = 8'd3;
    89: charMap = 8'd3;
    90: charMap = 8'd3;
    91: charMap = 8'd6;
    92: charMap = 8'd7;
    93: charMap = 8'd15;
    94: charMap = 8'd3;
    95: charMap = 8'd3;
    96: charMap = 8'd3;
    97: charMap = 8'd3;
    98: charMap = 8'd3;
    99: charMap = 8'd3;
    100: charMap = 8'd12;
    101: charMap = 8'd19;
    102: charMap = 8'd3;
    103: charMap = 8'd21;
    104: charMap = 8'd3;
    105: charMap = 8'd3;
    106: charMap = 8'd3;
    107: charMap = 8'd3;
    108: charMap = 8'd3;
    109: charMap = 8'd3;
    110: charMap = 8'd20;
    111: charMap = 8'd3;
    112: charMap = 8'd3;
    113: charMap = 8'd3;
    114: charMap = 8'd3;
    115: charMap = 8'd18;
    116: charMap = 8'd22;
    117: charMap = 8'd3;
    118: charMap = 8'd3;
    119: charMap = 8'd3;
    120: charMap = 8'd8;
    121: charMap = 8'd3;
    122: charMap = 8'd3;
    123: charMap = 8'd3;
    124: charMap = 8'd3;
    125: charMap = 8'd3;
    126: charMap = 8'd14;
    127: charMap = 8'd1;
    128: charMap = 8'd1;
    129: charMap = 8'd1;
    130: charMap = 8'd1;
    131: charMap = 8'd1;
    132: charMap = 8'd1;
    133: charMap = 8'd1;
    134: charMap = 8'd1;
    135: charMap = 8'd1;
    136: charMap = 8'd1;
    137: charMap = 8'd1;
    138: charMap = 8'd1;
    139: charMap = 8'd1;
    140: charMap = 8'd1;
    141: charMap = 8'd1;
    142: charMap = 8'd1;
    143: charMap = 8'd1;
    144: charMap = 8'd1;
    145: charMap = 8'd1;
    146: charMap = 8'd1;
    147: charMap = 8'd1;
    148: charMap = 8'd1;
    149: charMap = 8'd1;
    150: charMap = 8'd1;
    151: charMap = 8'd1;
    152: charMap = 8'd1;
    153: charMap = 8'd1;
    154: charMap = 8'd1;
    155: charMap = 8'd1;
    156: charMap = 8'd1;
    157: charMap = 8'd1;
    158: charMap = 8'd1;
    159: charMap = 8'd1;
    160: charMap = 8'd1;
    161: charMap = 8'd1;
    162: charMap = 8'd1;
    163: charMap = 8'd1;
    164: charMap = 8'd1;
    165: charMap = 8'd1;
    166: charMap = 8'd1;
    167: charMap = 8'd1;
    168: charMap = 8'd1;
    169: charMap = 8'd1;
    170: charMap = 8'd1;
    171: charMap = 8'd1;
    172: charMap = 8'd1;
    173: charMap = 8'd1;
    174: charMap = 8'd1;
    175: charMap = 8'd1;
    176: charMap = 8'd1;
    177: charMap = 8'd1;
    178: charMap = 8'd1;
    179: charMap = 8'd1;
    180: charMap = 8'd1;
    181: charMap = 8'd1;
    182: charMap = 8'd1;
    183: charMap = 8'd1;
    184: charMap = 8'd1;
    185: charMap = 8'd1;
    186: charMap = 8'd1;
    187: charMap = 8'd1;
    188: charMap = 8'd1;
    189: charMap = 8'd1;
    190: charMap = 8'd1;
    191: charMap = 8'd1;
    192: charMap = 8'd1;
    193: charMap = 8'd1;
    194: charMap = 8'd1;
    195: charMap = 8'd1;
    196: charMap = 8'd1;
    197: charMap = 8'd1;
    198: charMap = 8'd1;
    199: charMap = 8'd1;
    200: charMap = 8'd1;
    201: charMap = 8'd1;
    202: charMap = 8'd1;
    203: charMap = 8'd1;
    204: charMap = 8'd1;
    205: charMap = 8'd1;
    206: charMap = 8'd1;
    207: charMap = 8'd1;
    208: charMap = 8'd1;
    209: charMap = 8'd1;
    210: charMap = 8'd1;
    211: charMap = 8'd1;
    212: charMap = 8'd1;
    213: charMap = 8'd1;
    214: charMap = 8'd1;
    215: charMap = 8'd1;
    216: charMap = 8'd1;
    217: charMap = 8'd1;
    218: charMap = 8'd1;
    219: charMap = 8'd1;
    220: charMap = 8'd1;
    221: charMap = 8'd1;
    222: charMap = 8'd1;
    223: charMap = 8'd1;
    224: charMap = 8'd1;
    225: charMap = 8'd1;
    226: charMap = 8'd1;
    227: charMap = 8'd1;
    228: charMap = 8'd1;
    229: charMap = 8'd1;
    230: charMap = 8'd1;
    231: charMap = 8'd1;
    232: charMap = 8'd1;
    233: charMap = 8'd1;
    234: charMap = 8'd1;
    235: charMap = 8'd1;
    236: charMap = 8'd1;
    237: charMap = 8'd1;
    238: charMap = 8'd1;
    239: charMap = 8'd1;
    240: charMap = 8'd1;
    241: charMap = 8'd1;
    242: charMap = 8'd1;
    243: charMap = 8'd1;
    244: charMap = 8'd1;
    245: charMap = 8'd1;
    246: charMap = 8'd1;
    247: charMap = 8'd1;
    248: charMap = 8'd1;
    249: charMap = 8'd1;
    250: charMap = 8'd1;
    251: charMap = 8'd1;
    252: charMap = 8'd1;
    253: charMap = 8'd1;
    254: charMap = 8'd1;
    255: charMap = 8'd1;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd1;
    3: stateMap = 11'd2;
    4: stateMap = 11'd3;
    5: stateMap = 11'd4;
    6: stateMap = 11'd5;
    7: stateMap = 11'd6;
    8: stateMap = 11'd7;
    9: stateMap = 11'd8;
    10: stateMap = 11'd9;
    11: stateMap = 11'd10;
    12: stateMap = 11'd11;
    13: stateMap = 11'd12;
    14: stateMap = 11'd13;
    15: stateMap = 11'd14;
    16: stateMap = 11'd15;
    17: stateMap = 11'd16;
    18: stateMap = 11'd17;
    19: stateMap = 11'd18;
    20: stateMap = 11'd19;
    21: stateMap = 11'd20;
    22: stateMap = 11'd21;
    23: stateMap = 11'd22;
    24: stateMap = 11'd23;
    25: stateMap = 11'd24;
    26: stateMap = 11'd25;
    27: stateMap = 11'd26;
    28: stateMap = 11'd27;
    29: stateMap = 11'd28;
    30: stateMap = 11'd29;
    31: stateMap = 11'd30;
    32: stateMap = 11'd31;
    33: stateMap = 11'd32;
    34: stateMap = 11'd33;
    35: stateMap = 11'd34;
    36: stateMap = 11'd35;
    37: stateMap = 11'd36;
    38: stateMap = 11'd37;
    39: stateMap = 11'd38;
    40: stateMap = 11'd39;
    41: stateMap = 11'd40;
    42: stateMap = 11'd41;
    43: stateMap = 11'd42;
    44: stateMap = 11'd43;
    45: stateMap = 11'd44;
    46: stateMap = 11'd45;
    47: stateMap = 11'd46;
    48: stateMap = 11'd47;
    49: stateMap = 11'd48;
    50: stateMap = 11'd49;
    51: stateMap = 11'd50;
    52: stateMap = 11'd51;
    53: stateMap = 11'd52;
    54: stateMap = 11'd53;
    55: stateMap = 11'd54;
    56: stateMap = 11'd55;
    57: stateMap = 11'd56;
    58: stateMap = 11'd57;
    59: stateMap = 11'd13;
    60: stateMap = 11'd58;
    61: stateMap = 11'd59;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b1;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b0;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b0;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b0;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b0;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b0;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b0;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b0;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b0;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b0;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b0;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b0;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd3;
      3: stateTransition = 11'd3;
      4: stateTransition = 11'd3;
      5: stateTransition = 11'd3;
      6: stateTransition = 11'd3;
      7: stateTransition = 11'd3;
      8: stateTransition = 11'd3;
      9: stateTransition = 11'd3;
      10: stateTransition = 11'd3;
      11: stateTransition = 11'd3;
      12: stateTransition = 11'd3;
      13: stateTransition = 11'd3;
      14: stateTransition = 11'd3;
      15: stateTransition = 11'd3;
      16: stateTransition = 11'd3;
      17: stateTransition = 11'd5;
      18: stateTransition = 11'd3;
      19: stateTransition = 11'd3;
      20: stateTransition = 11'd3;
      21: stateTransition = 11'd3;
      22: stateTransition = 11'd3;
      23: stateTransition = 11'd1;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd6;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd2;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd6;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd7;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd56;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd8;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd8;
      6: stateTransition = 11'd8;
      7: stateTransition = 11'd8;
      8: stateTransition = 11'd8;
      9: stateTransition = 11'd8;
      10: stateTransition = 11'd8;
      11: stateTransition = 11'd8;
      12: stateTransition = 11'd8;
      13: stateTransition = 11'd8;
      14: stateTransition = 11'd8;
      15: stateTransition = 11'd8;
      16: stateTransition = 11'd8;
      17: stateTransition = 11'd8;
      18: stateTransition = 11'd8;
      19: stateTransition = 11'd8;
      20: stateTransition = 11'd8;
      21: stateTransition = 11'd8;
      22: stateTransition = 11'd8;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd9;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd8;
      4: stateTransition = 11'd11;
      5: stateTransition = 11'd8;
      6: stateTransition = 11'd8;
      7: stateTransition = 11'd8;
      8: stateTransition = 11'd8;
      9: stateTransition = 11'd8;
      10: stateTransition = 11'd8;
      11: stateTransition = 11'd8;
      12: stateTransition = 11'd8;
      13: stateTransition = 11'd8;
      14: stateTransition = 11'd8;
      15: stateTransition = 11'd8;
      16: stateTransition = 11'd8;
      17: stateTransition = 11'd8;
      18: stateTransition = 11'd8;
      19: stateTransition = 11'd8;
      20: stateTransition = 11'd8;
      21: stateTransition = 11'd8;
      22: stateTransition = 11'd8;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd12;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd13;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd14;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd15;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd13;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd57;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd57;
      6: stateTransition = 11'd57;
      7: stateTransition = 11'd57;
      8: stateTransition = 11'd57;
      9: stateTransition = 11'd57;
      10: stateTransition = 11'd57;
      11: stateTransition = 11'd57;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd57;
      14: stateTransition = 11'd57;
      15: stateTransition = 11'd57;
      16: stateTransition = 11'd57;
      17: stateTransition = 11'd57;
      18: stateTransition = 11'd57;
      19: stateTransition = 11'd57;
      20: stateTransition = 11'd57;
      21: stateTransition = 11'd57;
      22: stateTransition = 11'd57;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd17;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd17;
      10: stateTransition = 11'd17;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd17;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd17;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd18;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd61;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd20;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd21;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd22;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd23;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd25;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd28;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd29;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd30;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd31;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd32;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd33;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd34;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd35;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd36;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd37;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd38;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd39;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd40;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd41;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd42;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd43;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd44;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd45;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd46;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd47;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd48;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd49;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd51;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd52;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd2;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd54;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd55;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd2;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd2;
      10: stateTransition = 11'd2;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd2;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd4;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd10;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd57;
      4: stateTransition = 11'd16;
      5: stateTransition = 11'd57;
      6: stateTransition = 11'd57;
      7: stateTransition = 11'd57;
      8: stateTransition = 11'd57;
      9: stateTransition = 11'd57;
      10: stateTransition = 11'd57;
      11: stateTransition = 11'd57;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd57;
      14: stateTransition = 11'd57;
      15: stateTransition = 11'd57;
      16: stateTransition = 11'd57;
      17: stateTransition = 11'd57;
      18: stateTransition = 11'd57;
      19: stateTransition = 11'd57;
      20: stateTransition = 11'd57;
      21: stateTransition = 11'd57;
      22: stateTransition = 11'd57;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd26;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd26;
      10: stateTransition = 11'd26;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd26;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd26;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd58;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd58;
      10: stateTransition = 11'd58;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd58;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd58;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd60;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd60;
      10: stateTransition = 11'd60;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd60;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd60;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
