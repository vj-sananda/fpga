`define f0_W0_LSB  0
`define f0_W0_MSB  4

`define f1_W0_LSB  5
`define f1_W0_MSB  10

`define f2_W0_LSB  11
`define f2_W0_MSB  31
`define f2_W1_LSB  0
`define f2_W1_MSB  10

`define f3_W1_LSB  11
`define f3_W1_MSB  31
`define f3_W2_LSB  0
`define f3_W2_MSB  8

`define f4_W2_LSB  9
`define f4_W2_MSB  31

