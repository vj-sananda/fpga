   //Define bitvector widths
   parameter w_din = 32,
	       w_f0 = 5,
	       w_f1 = 6,
	       w_f2 = 32,
	       w_f3 = 30,
	       w_f4 = 23;

   parameter msb_states=2;//Num states 
