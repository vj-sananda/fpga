`timescale 1ns/1ps

`define ENABLED_REGEX_CATEGORY_dhcp TRUE

module CATEGORY_dhcp_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_CATEGORY_dhcp

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd4;
    1: charMap = 8'd1;
    2: charMap = 8'd1;
    3: charMap = 8'd5;
    4: charMap = 8'd5;
    5: charMap = 8'd5;
    6: charMap = 8'd3;
    7: charMap = 8'd5;
    8: charMap = 8'd5;
    9: charMap = 8'd5;
    10: charMap = 8'd2;
    11: charMap = 8'd5;
    12: charMap = 8'd5;
    13: charMap = 8'd2;
    14: charMap = 8'd5;
    15: charMap = 8'd5;
    16: charMap = 8'd5;
    17: charMap = 8'd5;
    18: charMap = 8'd5;
    19: charMap = 8'd5;
    20: charMap = 8'd5;
    21: charMap = 8'd5;
    22: charMap = 8'd5;
    23: charMap = 8'd5;
    24: charMap = 8'd5;
    25: charMap = 8'd5;
    26: charMap = 8'd5;
    27: charMap = 8'd5;
    28: charMap = 8'd5;
    29: charMap = 8'd5;
    30: charMap = 8'd5;
    31: charMap = 8'd5;
    32: charMap = 8'd5;
    33: charMap = 8'd4;
    34: charMap = 8'd4;
    35: charMap = 8'd4;
    36: charMap = 8'd4;
    37: charMap = 8'd4;
    38: charMap = 8'd4;
    39: charMap = 8'd4;
    40: charMap = 8'd4;
    41: charMap = 8'd4;
    42: charMap = 8'd4;
    43: charMap = 8'd4;
    44: charMap = 8'd4;
    45: charMap = 8'd4;
    46: charMap = 8'd4;
    47: charMap = 8'd4;
    48: charMap = 8'd4;
    49: charMap = 8'd4;
    50: charMap = 8'd4;
    51: charMap = 8'd4;
    52: charMap = 8'd4;
    53: charMap = 8'd4;
    54: charMap = 8'd4;
    55: charMap = 8'd4;
    56: charMap = 8'd4;
    57: charMap = 8'd4;
    58: charMap = 8'd4;
    59: charMap = 8'd4;
    60: charMap = 8'd4;
    61: charMap = 8'd4;
    62: charMap = 8'd4;
    63: charMap = 8'd4;
    64: charMap = 8'd4;
    65: charMap = 8'd4;
    66: charMap = 8'd4;
    67: charMap = 8'd4;
    68: charMap = 8'd4;
    69: charMap = 8'd4;
    70: charMap = 8'd4;
    71: charMap = 8'd4;
    72: charMap = 8'd4;
    73: charMap = 8'd4;
    74: charMap = 8'd4;
    75: charMap = 8'd4;
    76: charMap = 8'd4;
    77: charMap = 8'd4;
    78: charMap = 8'd4;
    79: charMap = 8'd4;
    80: charMap = 8'd4;
    81: charMap = 8'd4;
    82: charMap = 8'd4;
    83: charMap = 8'd4;
    84: charMap = 8'd4;
    85: charMap = 8'd4;
    86: charMap = 8'd4;
    87: charMap = 8'd4;
    88: charMap = 8'd4;
    89: charMap = 8'd4;
    90: charMap = 8'd4;
    91: charMap = 8'd4;
    92: charMap = 8'd4;
    93: charMap = 8'd4;
    94: charMap = 8'd4;
    95: charMap = 8'd4;
    96: charMap = 8'd4;
    97: charMap = 8'd4;
    98: charMap = 8'd4;
    99: charMap = 8'd6;
    100: charMap = 8'd4;
    101: charMap = 8'd4;
    102: charMap = 8'd4;
    103: charMap = 8'd4;
    104: charMap = 8'd4;
    105: charMap = 8'd4;
    106: charMap = 8'd4;
    107: charMap = 8'd4;
    108: charMap = 8'd4;
    109: charMap = 8'd4;
    110: charMap = 8'd4;
    111: charMap = 8'd4;
    112: charMap = 8'd4;
    113: charMap = 8'd4;
    114: charMap = 8'd4;
    115: charMap = 8'd8;
    116: charMap = 8'd4;
    117: charMap = 8'd4;
    118: charMap = 8'd4;
    119: charMap = 8'd4;
    120: charMap = 8'd4;
    121: charMap = 8'd4;
    122: charMap = 8'd4;
    123: charMap = 8'd4;
    124: charMap = 8'd4;
    125: charMap = 8'd4;
    126: charMap = 8'd4;
    127: charMap = 8'd4;
    128: charMap = 8'd4;
    129: charMap = 8'd4;
    130: charMap = 8'd7;
    131: charMap = 8'd4;
    132: charMap = 8'd4;
    133: charMap = 8'd4;
    134: charMap = 8'd4;
    135: charMap = 8'd4;
    136: charMap = 8'd4;
    137: charMap = 8'd4;
    138: charMap = 8'd4;
    139: charMap = 8'd4;
    140: charMap = 8'd4;
    141: charMap = 8'd4;
    142: charMap = 8'd4;
    143: charMap = 8'd4;
    144: charMap = 8'd4;
    145: charMap = 8'd4;
    146: charMap = 8'd4;
    147: charMap = 8'd4;
    148: charMap = 8'd4;
    149: charMap = 8'd4;
    150: charMap = 8'd4;
    151: charMap = 8'd4;
    152: charMap = 8'd4;
    153: charMap = 8'd4;
    154: charMap = 8'd4;
    155: charMap = 8'd4;
    156: charMap = 8'd4;
    157: charMap = 8'd4;
    158: charMap = 8'd4;
    159: charMap = 8'd4;
    160: charMap = 8'd4;
    161: charMap = 8'd4;
    162: charMap = 8'd4;
    163: charMap = 8'd4;
    164: charMap = 8'd4;
    165: charMap = 8'd4;
    166: charMap = 8'd4;
    167: charMap = 8'd4;
    168: charMap = 8'd4;
    169: charMap = 8'd4;
    170: charMap = 8'd4;
    171: charMap = 8'd4;
    172: charMap = 8'd4;
    173: charMap = 8'd4;
    174: charMap = 8'd4;
    175: charMap = 8'd4;
    176: charMap = 8'd4;
    177: charMap = 8'd4;
    178: charMap = 8'd4;
    179: charMap = 8'd4;
    180: charMap = 8'd4;
    181: charMap = 8'd4;
    182: charMap = 8'd4;
    183: charMap = 8'd4;
    184: charMap = 8'd4;
    185: charMap = 8'd4;
    186: charMap = 8'd4;
    187: charMap = 8'd4;
    188: charMap = 8'd4;
    189: charMap = 8'd4;
    190: charMap = 8'd4;
    191: charMap = 8'd4;
    192: charMap = 8'd4;
    193: charMap = 8'd4;
    194: charMap = 8'd4;
    195: charMap = 8'd4;
    196: charMap = 8'd4;
    197: charMap = 8'd4;
    198: charMap = 8'd4;
    199: charMap = 8'd4;
    200: charMap = 8'd4;
    201: charMap = 8'd4;
    202: charMap = 8'd4;
    203: charMap = 8'd4;
    204: charMap = 8'd4;
    205: charMap = 8'd4;
    206: charMap = 8'd4;
    207: charMap = 8'd4;
    208: charMap = 8'd4;
    209: charMap = 8'd4;
    210: charMap = 8'd4;
    211: charMap = 8'd4;
    212: charMap = 8'd4;
    213: charMap = 8'd4;
    214: charMap = 8'd4;
    215: charMap = 8'd4;
    216: charMap = 8'd4;
    217: charMap = 8'd4;
    218: charMap = 8'd4;
    219: charMap = 8'd4;
    220: charMap = 8'd4;
    221: charMap = 8'd4;
    222: charMap = 8'd4;
    223: charMap = 8'd4;
    224: charMap = 8'd4;
    225: charMap = 8'd4;
    226: charMap = 8'd4;
    227: charMap = 8'd4;
    228: charMap = 8'd4;
    229: charMap = 8'd4;
    230: charMap = 8'd4;
    231: charMap = 8'd4;
    232: charMap = 8'd4;
    233: charMap = 8'd4;
    234: charMap = 8'd4;
    235: charMap = 8'd4;
    236: charMap = 8'd4;
    237: charMap = 8'd4;
    238: charMap = 8'd4;
    239: charMap = 8'd4;
    240: charMap = 8'd4;
    241: charMap = 8'd4;
    242: charMap = 8'd4;
    243: charMap = 8'd4;
    244: charMap = 8'd4;
    245: charMap = 8'd4;
    246: charMap = 8'd4;
    247: charMap = 8'd4;
    248: charMap = 8'd4;
    249: charMap = 8'd4;
    250: charMap = 8'd4;
    251: charMap = 8'd4;
    252: charMap = 8'd4;
    253: charMap = 8'd4;
    254: charMap = 8'd4;
    255: charMap = 8'd4;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd2;
    3: stateMap = 11'd3;
    4: stateMap = 11'd4;
    5: stateMap = 11'd5;
    6: stateMap = 11'd6;
    7: stateMap = 11'd7;
    8: stateMap = 11'd2;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b0;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b0;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd1;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd5;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd5;
      5: stateTransition = 11'd5;
      6: stateTransition = 11'd8;
      7: stateTransition = 11'd7;
      8: stateTransition = 11'd5;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd4;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd4;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd4;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd5;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd5;
      5: stateTransition = 11'd5;
      6: stateTransition = 11'd8;
      7: stateTransition = 11'd5;
      8: stateTransition = 11'd5;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd5;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd5;
      5: stateTransition = 11'd5;
      6: stateTransition = 11'd2;
      7: stateTransition = 11'd5;
      8: stateTransition = 11'd5;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd5;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd5;
      5: stateTransition = 11'd5;
      6: stateTransition = 11'd8;
      7: stateTransition = 11'd5;
      8: stateTransition = 11'd6;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
