`include "pkt.defn.vh"

`define F0_W 5
`define F1_W 6
`define F2_W 32
`define F3_W 30
`define F4_W 23

