`timescale 1ns/1ps

`define ENABLED_REGEX_CATEGORY_fasttrack TRUE

module CATEGORY_fasttrack_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_CATEGORY_fasttrack

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd6;
    1: charMap = 8'd6;
    2: charMap = 8'd6;
    3: charMap = 8'd6;
    4: charMap = 8'd6;
    5: charMap = 8'd6;
    6: charMap = 8'd6;
    7: charMap = 8'd6;
    8: charMap = 8'd6;
    9: charMap = 8'd6;
    10: charMap = 8'd0;
    11: charMap = 8'd6;
    12: charMap = 8'd6;
    13: charMap = 8'd0;
    14: charMap = 8'd6;
    15: charMap = 8'd6;
    16: charMap = 8'd6;
    17: charMap = 8'd6;
    18: charMap = 8'd6;
    19: charMap = 8'd6;
    20: charMap = 8'd6;
    21: charMap = 8'd6;
    22: charMap = 8'd6;
    23: charMap = 8'd6;
    24: charMap = 8'd6;
    25: charMap = 8'd6;
    26: charMap = 8'd6;
    27: charMap = 8'd6;
    28: charMap = 8'd6;
    29: charMap = 8'd6;
    30: charMap = 8'd6;
    31: charMap = 8'd6;
    32: charMap = 8'd4;
    33: charMap = 8'd13;
    34: charMap = 8'd13;
    35: charMap = 8'd13;
    36: charMap = 8'd13;
    37: charMap = 8'd13;
    38: charMap = 8'd13;
    39: charMap = 8'd13;
    40: charMap = 8'd13;
    41: charMap = 8'd13;
    42: charMap = 8'd13;
    43: charMap = 8'd13;
    44: charMap = 8'd13;
    45: charMap = 8'd25;
    46: charMap = 8'd13;
    47: charMap = 8'd5;
    48: charMap = 8'd31;
    49: charMap = 8'd24;
    50: charMap = 8'd31;
    51: charMap = 8'd31;
    52: charMap = 8'd31;
    53: charMap = 8'd31;
    54: charMap = 8'd31;
    55: charMap = 8'd31;
    56: charMap = 8'd31;
    57: charMap = 8'd31;
    58: charMap = 8'd26;
    59: charMap = 8'd13;
    60: charMap = 8'd13;
    61: charMap = 8'd22;
    62: charMap = 8'd13;
    63: charMap = 8'd13;
    64: charMap = 8'd13;
    65: charMap = 8'd13;
    66: charMap = 8'd13;
    67: charMap = 8'd13;
    68: charMap = 8'd13;
    69: charMap = 8'd13;
    70: charMap = 8'd13;
    71: charMap = 8'd13;
    72: charMap = 8'd13;
    73: charMap = 8'd13;
    74: charMap = 8'd13;
    75: charMap = 8'd13;
    76: charMap = 8'd13;
    77: charMap = 8'd13;
    78: charMap = 8'd13;
    79: charMap = 8'd13;
    80: charMap = 8'd13;
    81: charMap = 8'd13;
    82: charMap = 8'd13;
    83: charMap = 8'd13;
    84: charMap = 8'd13;
    85: charMap = 8'd13;
    86: charMap = 8'd13;
    87: charMap = 8'd13;
    88: charMap = 8'd13;
    89: charMap = 8'd13;
    90: charMap = 8'd13;
    91: charMap = 8'd13;
    92: charMap = 8'd13;
    93: charMap = 8'd13;
    94: charMap = 8'd13;
    95: charMap = 8'd13;
    96: charMap = 8'd13;
    97: charMap = 8'd12;
    98: charMap = 8'd23;
    99: charMap = 8'd23;
    100: charMap = 8'd7;
    101: charMap = 8'd2;
    102: charMap = 8'd19;
    103: charMap = 8'd1;
    104: charMap = 8'd21;
    105: charMap = 8'd20;
    106: charMap = 8'd13;
    107: charMap = 8'd18;
    108: charMap = 8'd11;
    109: charMap = 8'd29;
    110: charMap = 8'd10;
    111: charMap = 8'd8;
    112: charMap = 8'd16;
    113: charMap = 8'd13;
    114: charMap = 8'd17;
    115: charMap = 8'd14;
    116: charMap = 8'd3;
    117: charMap = 8'd15;
    118: charMap = 8'd30;
    119: charMap = 8'd9;
    120: charMap = 8'd28;
    121: charMap = 8'd13;
    122: charMap = 8'd27;
    123: charMap = 8'd13;
    124: charMap = 8'd13;
    125: charMap = 8'd13;
    126: charMap = 8'd13;
    127: charMap = 8'd6;
    128: charMap = 8'd6;
    129: charMap = 8'd6;
    130: charMap = 8'd6;
    131: charMap = 8'd6;
    132: charMap = 8'd6;
    133: charMap = 8'd6;
    134: charMap = 8'd6;
    135: charMap = 8'd6;
    136: charMap = 8'd6;
    137: charMap = 8'd6;
    138: charMap = 8'd6;
    139: charMap = 8'd6;
    140: charMap = 8'd6;
    141: charMap = 8'd6;
    142: charMap = 8'd6;
    143: charMap = 8'd6;
    144: charMap = 8'd6;
    145: charMap = 8'd6;
    146: charMap = 8'd6;
    147: charMap = 8'd6;
    148: charMap = 8'd6;
    149: charMap = 8'd6;
    150: charMap = 8'd6;
    151: charMap = 8'd6;
    152: charMap = 8'd6;
    153: charMap = 8'd6;
    154: charMap = 8'd6;
    155: charMap = 8'd6;
    156: charMap = 8'd6;
    157: charMap = 8'd6;
    158: charMap = 8'd6;
    159: charMap = 8'd6;
    160: charMap = 8'd6;
    161: charMap = 8'd6;
    162: charMap = 8'd6;
    163: charMap = 8'd6;
    164: charMap = 8'd6;
    165: charMap = 8'd6;
    166: charMap = 8'd6;
    167: charMap = 8'd6;
    168: charMap = 8'd6;
    169: charMap = 8'd6;
    170: charMap = 8'd6;
    171: charMap = 8'd6;
    172: charMap = 8'd6;
    173: charMap = 8'd6;
    174: charMap = 8'd6;
    175: charMap = 8'd6;
    176: charMap = 8'd6;
    177: charMap = 8'd6;
    178: charMap = 8'd6;
    179: charMap = 8'd6;
    180: charMap = 8'd6;
    181: charMap = 8'd6;
    182: charMap = 8'd6;
    183: charMap = 8'd6;
    184: charMap = 8'd6;
    185: charMap = 8'd6;
    186: charMap = 8'd6;
    187: charMap = 8'd6;
    188: charMap = 8'd6;
    189: charMap = 8'd6;
    190: charMap = 8'd6;
    191: charMap = 8'd6;
    192: charMap = 8'd6;
    193: charMap = 8'd6;
    194: charMap = 8'd6;
    195: charMap = 8'd6;
    196: charMap = 8'd6;
    197: charMap = 8'd6;
    198: charMap = 8'd6;
    199: charMap = 8'd6;
    200: charMap = 8'd6;
    201: charMap = 8'd6;
    202: charMap = 8'd6;
    203: charMap = 8'd6;
    204: charMap = 8'd6;
    205: charMap = 8'd6;
    206: charMap = 8'd6;
    207: charMap = 8'd6;
    208: charMap = 8'd6;
    209: charMap = 8'd6;
    210: charMap = 8'd6;
    211: charMap = 8'd6;
    212: charMap = 8'd6;
    213: charMap = 8'd6;
    214: charMap = 8'd6;
    215: charMap = 8'd6;
    216: charMap = 8'd6;
    217: charMap = 8'd6;
    218: charMap = 8'd6;
    219: charMap = 8'd6;
    220: charMap = 8'd6;
    221: charMap = 8'd6;
    222: charMap = 8'd6;
    223: charMap = 8'd6;
    224: charMap = 8'd6;
    225: charMap = 8'd6;
    226: charMap = 8'd6;
    227: charMap = 8'd6;
    228: charMap = 8'd6;
    229: charMap = 8'd6;
    230: charMap = 8'd6;
    231: charMap = 8'd6;
    232: charMap = 8'd6;
    233: charMap = 8'd6;
    234: charMap = 8'd6;
    235: charMap = 8'd6;
    236: charMap = 8'd6;
    237: charMap = 8'd6;
    238: charMap = 8'd6;
    239: charMap = 8'd6;
    240: charMap = 8'd6;
    241: charMap = 8'd6;
    242: charMap = 8'd6;
    243: charMap = 8'd6;
    244: charMap = 8'd6;
    245: charMap = 8'd6;
    246: charMap = 8'd6;
    247: charMap = 8'd6;
    248: charMap = 8'd6;
    249: charMap = 8'd6;
    250: charMap = 8'd6;
    251: charMap = 8'd6;
    252: charMap = 8'd6;
    253: charMap = 8'd6;
    254: charMap = 8'd6;
    255: charMap = 8'd6;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd1;
    3: stateMap = 11'd2;
    4: stateMap = 11'd3;
    5: stateMap = 11'd4;
    6: stateMap = 11'd5;
    7: stateMap = 11'd6;
    8: stateMap = 11'd7;
    9: stateMap = 11'd8;
    10: stateMap = 11'd9;
    11: stateMap = 11'd10;
    12: stateMap = 11'd11;
    13: stateMap = 11'd12;
    14: stateMap = 11'd13;
    15: stateMap = 11'd14;
    16: stateMap = 11'd15;
    17: stateMap = 11'd16;
    18: stateMap = 11'd17;
    19: stateMap = 11'd18;
    20: stateMap = 11'd19;
    21: stateMap = 11'd20;
    22: stateMap = 11'd21;
    23: stateMap = 11'd22;
    24: stateMap = 11'd23;
    25: stateMap = 11'd24;
    26: stateMap = 11'd25;
    27: stateMap = 11'd26;
    28: stateMap = 11'd27;
    29: stateMap = 11'd28;
    30: stateMap = 11'd29;
    31: stateMap = 11'd30;
    32: stateMap = 11'd31;
    33: stateMap = 11'd32;
    34: stateMap = 11'd33;
    35: stateMap = 11'd34;
    36: stateMap = 11'd35;
    37: stateMap = 11'd36;
    38: stateMap = 11'd37;
    39: stateMap = 11'd38;
    40: stateMap = 11'd39;
    41: stateMap = 11'd40;
    42: stateMap = 11'd41;
    43: stateMap = 11'd42;
    44: stateMap = 11'd43;
    45: stateMap = 11'd44;
    46: stateMap = 11'd45;
    47: stateMap = 11'd46;
    48: stateMap = 11'd47;
    49: stateMap = 11'd48;
    50: stateMap = 11'd49;
    51: stateMap = 11'd50;
    52: stateMap = 11'd51;
    53: stateMap = 11'd52;
    54: stateMap = 11'd53;
    55: stateMap = 11'd54;
    56: stateMap = 11'd55;
    57: stateMap = 11'd56;
    58: stateMap = 11'd57;
    59: stateMap = 11'd58;
    60: stateMap = 11'd59;
    61: stateMap = 11'd60;
    62: stateMap = 11'd61;
    63: stateMap = 11'd62;
    64: stateMap = 11'd63;
    65: stateMap = 11'd64;
    66: stateMap = 11'd65;
    67: stateMap = 11'd66;
    68: stateMap = 11'd7;
    69: stateMap = 11'd67;
    70: stateMap = 11'd68;
    71: stateMap = 11'd69;
    72: stateMap = 11'd70;
    73: stateMap = 11'd71;
    74: stateMap = 11'd72;
    75: stateMap = 11'd73;
    76: stateMap = 11'd74;
    77: stateMap = 11'd75;
    78: stateMap = 11'd76;
    79: stateMap = 11'd77;
    80: stateMap = 11'd78;
    81: stateMap = 11'd79;
    82: stateMap = 11'd80;
    83: stateMap = 11'd81;
    84: stateMap = 11'd82;
    85: stateMap = 11'd83;
    86: stateMap = 11'd84;
    87: stateMap = 11'd85;
    88: stateMap = 11'd86;
    89: stateMap = 11'd87;
    90: stateMap = 11'd88;
    91: stateMap = 11'd89;
    92: stateMap = 11'd90;
    93: stateMap = 11'd91;
    94: stateMap = 11'd92;
    95: stateMap = 11'd93;
    96: stateMap = 11'd94;
    97: stateMap = 11'd95;
    98: stateMap = 11'd96;
    99: stateMap = 11'd57;
    100: stateMap = 11'd97;
    101: stateMap = 11'd98;
    102: stateMap = 11'd99;
    103: stateMap = 11'd100;
    104: stateMap = 11'd101;
    105: stateMap = 11'd102;
    106: stateMap = 11'd103;
    107: stateMap = 11'd104;
    108: stateMap = 11'd105;
    109: stateMap = 11'd106;
    110: stateMap = 11'd107;
    111: stateMap = 11'd108;
    112: stateMap = 11'd109;
    113: stateMap = 11'd110;
    114: stateMap = 11'd111;
    115: stateMap = 11'd112;
    116: stateMap = 11'd113;
    117: stateMap = 11'd114;
    118: stateMap = 11'd115;
    119: stateMap = 11'd116;
    120: stateMap = 11'd117;
    121: stateMap = 11'd118;
    122: stateMap = 11'd119;
    123: stateMap = 11'd120;
    124: stateMap = 11'd121;
    125: stateMap = 11'd122;
    126: stateMap = 11'd123;
    127: stateMap = 11'd124;
    128: stateMap = 11'd125;
    129: stateMap = 11'd126;
    130: stateMap = 11'd127;
    131: stateMap = 11'd128;
    132: stateMap = 11'd129;
    133: stateMap = 11'd130;
    134: stateMap = 11'd131;
    135: stateMap = 11'd132;
    136: stateMap = 11'd133;
    137: stateMap = 11'd134;
    138: stateMap = 11'd135;
    139: stateMap = 11'd136;
    140: stateMap = 11'd137;
    141: stateMap = 11'd138;
    142: stateMap = 11'd139;
    143: stateMap = 11'd140;
    144: stateMap = 11'd141;
    145: stateMap = 11'd142;
    146: stateMap = 11'd143;
    147: stateMap = 11'd144;
    148: stateMap = 11'd145;
    149: stateMap = 11'd146;
    150: stateMap = 11'd147;
    151: stateMap = 11'd148;
    152: stateMap = 11'd145;
    153: stateMap = 11'd145;
    154: stateMap = 11'd149;
    155: stateMap = 11'd150;
    156: stateMap = 11'd147;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b1;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b1;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b1;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b0;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b0;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b0;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b0;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b0;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b0;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b0;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b0;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b0;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b0;
    62: acceptStates = 1'b0;
    63: acceptStates = 1'b0;
    64: acceptStates = 1'b0;
    65: acceptStates = 1'b0;
    66: acceptStates = 1'b0;
    67: acceptStates = 1'b0;
    68: acceptStates = 1'b0;
    69: acceptStates = 1'b0;
    70: acceptStates = 1'b0;
    71: acceptStates = 1'b0;
    72: acceptStates = 1'b0;
    73: acceptStates = 1'b0;
    74: acceptStates = 1'b0;
    75: acceptStates = 1'b0;
    76: acceptStates = 1'b0;
    77: acceptStates = 1'b0;
    78: acceptStates = 1'b0;
    79: acceptStates = 1'b0;
    80: acceptStates = 1'b0;
    81: acceptStates = 1'b0;
    82: acceptStates = 1'b0;
    83: acceptStates = 1'b0;
    84: acceptStates = 1'b0;
    85: acceptStates = 1'b0;
    86: acceptStates = 1'b0;
    87: acceptStates = 1'b0;
    88: acceptStates = 1'b0;
    89: acceptStates = 1'b0;
    90: acceptStates = 1'b0;
    91: acceptStates = 1'b0;
    92: acceptStates = 1'b0;
    93: acceptStates = 1'b0;
    94: acceptStates = 1'b0;
    95: acceptStates = 1'b0;
    96: acceptStates = 1'b0;
    97: acceptStates = 1'b1;
    98: acceptStates = 1'b0;
    99: acceptStates = 1'b0;
    100: acceptStates = 1'b0;
    101: acceptStates = 1'b0;
    102: acceptStates = 1'b0;
    103: acceptStates = 1'b0;
    104: acceptStates = 1'b0;
    105: acceptStates = 1'b0;
    106: acceptStates = 1'b0;
    107: acceptStates = 1'b0;
    108: acceptStates = 1'b0;
    109: acceptStates = 1'b0;
    110: acceptStates = 1'b0;
    111: acceptStates = 1'b0;
    112: acceptStates = 1'b0;
    113: acceptStates = 1'b0;
    114: acceptStates = 1'b0;
    115: acceptStates = 1'b0;
    116: acceptStates = 1'b0;
    117: acceptStates = 1'b0;
    118: acceptStates = 1'b0;
    119: acceptStates = 1'b0;
    120: acceptStates = 1'b0;
    121: acceptStates = 1'b0;
    122: acceptStates = 1'b0;
    123: acceptStates = 1'b0;
    124: acceptStates = 1'b0;
    125: acceptStates = 1'b0;
    126: acceptStates = 1'b0;
    127: acceptStates = 1'b0;
    128: acceptStates = 1'b0;
    129: acceptStates = 1'b0;
    130: acceptStates = 1'b0;
    131: acceptStates = 1'b0;
    132: acceptStates = 1'b0;
    133: acceptStates = 1'b0;
    134: acceptStates = 1'b0;
    135: acceptStates = 1'b0;
    136: acceptStates = 1'b0;
    137: acceptStates = 1'b0;
    138: acceptStates = 1'b0;
    139: acceptStates = 1'b0;
    140: acceptStates = 1'b0;
    141: acceptStates = 1'b0;
    142: acceptStates = 1'b0;
    143: acceptStates = 1'b0;
    144: acceptStates = 1'b0;
    145: acceptStates = 1'b0;
    146: acceptStates = 1'b0;
    147: acceptStates = 1'b0;
    148: acceptStates = 1'b0;
    149: acceptStates = 1'b0;
    150: acceptStates = 1'b0;
    151: acceptStates = 1'b0;
    152: acceptStates = 1'b1;
    153: acceptStates = 1'b0;
    154: acceptStates = 1'b0;
    155: acceptStates = 1'b0;
    156: acceptStates = 1'b1;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd5;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd7;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd1;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd9;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd10;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd97;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd97;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd2;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd2;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd12;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd68;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd98;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd14;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd15;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd16;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd18;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd20;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd21;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd22;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd101;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd23;
      2: stateTransition = 11'd23;
      3: stateTransition = 11'd23;
      4: stateTransition = 11'd23;
      5: stateTransition = 11'd23;
      6: stateTransition = 11'd23;
      7: stateTransition = 11'd23;
      8: stateTransition = 11'd23;
      9: stateTransition = 11'd23;
      10: stateTransition = 11'd23;
      11: stateTransition = 11'd23;
      12: stateTransition = 11'd23;
      13: stateTransition = 11'd23;
      14: stateTransition = 11'd23;
      15: stateTransition = 11'd23;
      16: stateTransition = 11'd23;
      17: stateTransition = 11'd23;
      18: stateTransition = 11'd23;
      19: stateTransition = 11'd23;
      20: stateTransition = 11'd23;
      21: stateTransition = 11'd23;
      22: stateTransition = 11'd23;
      23: stateTransition = 11'd23;
      24: stateTransition = 11'd23;
      25: stateTransition = 11'd23;
      26: stateTransition = 11'd23;
      27: stateTransition = 11'd23;
      28: stateTransition = 11'd23;
      29: stateTransition = 11'd23;
      30: stateTransition = 11'd23;
      31: stateTransition = 11'd23;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd135;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd135;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd26;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd28;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd29;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd102;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd103;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd30;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd31;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd32;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd33;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd34;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd35;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd104;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd38;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd39;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd40;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd41;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd107;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd42;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd106;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd121;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd44;
      15: stateTransition = 11'd45;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd46;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd47;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd49;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd108;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd50;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd51;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd2;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd54;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd55;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd2;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd124;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd110;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd111;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd57;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd112;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd61;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd129;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd62;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd65;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd66;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd67;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd59;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd4;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd4;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    60: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd115;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    61: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd69;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    62: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd71;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    63: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd153;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    64: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd99;
      2: stateTransition = 11'd99;
      3: stateTransition = 11'd99;
      4: stateTransition = 11'd99;
      5: stateTransition = 11'd99;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd99;
      8: stateTransition = 11'd99;
      9: stateTransition = 11'd99;
      10: stateTransition = 11'd99;
      11: stateTransition = 11'd99;
      12: stateTransition = 11'd99;
      13: stateTransition = 11'd99;
      14: stateTransition = 11'd99;
      15: stateTransition = 11'd99;
      16: stateTransition = 11'd99;
      17: stateTransition = 11'd99;
      18: stateTransition = 11'd99;
      19: stateTransition = 11'd99;
      20: stateTransition = 11'd99;
      21: stateTransition = 11'd99;
      22: stateTransition = 11'd99;
      23: stateTransition = 11'd99;
      24: stateTransition = 11'd99;
      25: stateTransition = 11'd99;
      26: stateTransition = 11'd99;
      27: stateTransition = 11'd99;
      28: stateTransition = 11'd99;
      29: stateTransition = 11'd99;
      30: stateTransition = 11'd99;
      31: stateTransition = 11'd99;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    65: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd118;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    66: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd72;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    67: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd120;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    68: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd75;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd76;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    69: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd77;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    70: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd119;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    71: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd79;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    72: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd80;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    73: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd76;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    74: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd2;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    75: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    76: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd65;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    77: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd84;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    78: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd2;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    79: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd85;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    80: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd86;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    81: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd87;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    82: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd88;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    83: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd89;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    84: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd2;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    85: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd90;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    86: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd2;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    87: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd91;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    88: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd92;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    89: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd46;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    90: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd93;
      2: stateTransition = 11'd93;
      3: stateTransition = 11'd93;
      4: stateTransition = 11'd93;
      5: stateTransition = 11'd93;
      6: stateTransition = 11'd93;
      7: stateTransition = 11'd93;
      8: stateTransition = 11'd93;
      9: stateTransition = 11'd93;
      10: stateTransition = 11'd93;
      11: stateTransition = 11'd93;
      12: stateTransition = 11'd93;
      13: stateTransition = 11'd93;
      14: stateTransition = 11'd93;
      15: stateTransition = 11'd93;
      16: stateTransition = 11'd93;
      17: stateTransition = 11'd93;
      18: stateTransition = 11'd93;
      19: stateTransition = 11'd93;
      20: stateTransition = 11'd93;
      21: stateTransition = 11'd93;
      22: stateTransition = 11'd93;
      23: stateTransition = 11'd93;
      24: stateTransition = 11'd93;
      25: stateTransition = 11'd93;
      26: stateTransition = 11'd93;
      27: stateTransition = 11'd93;
      28: stateTransition = 11'd93;
      29: stateTransition = 11'd93;
      30: stateTransition = 11'd93;
      31: stateTransition = 11'd93;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    91: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd2;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    92: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd95;
      2: stateTransition = 11'd95;
      3: stateTransition = 11'd95;
      4: stateTransition = 11'd137;
      5: stateTransition = 11'd95;
      6: stateTransition = 11'd93;
      7: stateTransition = 11'd95;
      8: stateTransition = 11'd95;
      9: stateTransition = 11'd95;
      10: stateTransition = 11'd95;
      11: stateTransition = 11'd95;
      12: stateTransition = 11'd95;
      13: stateTransition = 11'd95;
      14: stateTransition = 11'd95;
      15: stateTransition = 11'd95;
      16: stateTransition = 11'd95;
      17: stateTransition = 11'd95;
      18: stateTransition = 11'd95;
      19: stateTransition = 11'd95;
      20: stateTransition = 11'd95;
      21: stateTransition = 11'd95;
      22: stateTransition = 11'd95;
      23: stateTransition = 11'd95;
      24: stateTransition = 11'd95;
      25: stateTransition = 11'd95;
      26: stateTransition = 11'd95;
      27: stateTransition = 11'd95;
      28: stateTransition = 11'd95;
      29: stateTransition = 11'd95;
      30: stateTransition = 11'd95;
      31: stateTransition = 11'd95;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    93: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd8;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    94: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd155;
      2: stateTransition = 11'd155;
      3: stateTransition = 11'd155;
      4: stateTransition = 11'd139;
      5: stateTransition = 11'd155;
      6: stateTransition = 11'd93;
      7: stateTransition = 11'd155;
      8: stateTransition = 11'd155;
      9: stateTransition = 11'd155;
      10: stateTransition = 11'd155;
      11: stateTransition = 11'd155;
      12: stateTransition = 11'd155;
      13: stateTransition = 11'd155;
      14: stateTransition = 11'd155;
      15: stateTransition = 11'd155;
      16: stateTransition = 11'd155;
      17: stateTransition = 11'd155;
      18: stateTransition = 11'd155;
      19: stateTransition = 11'd155;
      20: stateTransition = 11'd155;
      21: stateTransition = 11'd155;
      22: stateTransition = 11'd155;
      23: stateTransition = 11'd155;
      24: stateTransition = 11'd155;
      25: stateTransition = 11'd155;
      26: stateTransition = 11'd155;
      27: stateTransition = 11'd155;
      28: stateTransition = 11'd155;
      29: stateTransition = 11'd155;
      30: stateTransition = 11'd155;
      31: stateTransition = 11'd155;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    95: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd6;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd6;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    96: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd17;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    97: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd60;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd60;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    98: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd25;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    99: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd36;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    100: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    101: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd43;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    102: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd48;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    103: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd52;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    104: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd109;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    105: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd56;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    106: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd58;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    107: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd63;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    108: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    109: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd114;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    110: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd70;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    111: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    112: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd74;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    113: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd94;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    114: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd81;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    115: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd78;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    116: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd83;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    117: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd82;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    118: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    119: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd96;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    120: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd100;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd100;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    121: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd113;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    122: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd117;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    123: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd116;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd68;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    124: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd122;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd150;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    125: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd123;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd123;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    126: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd125;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    127: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd68;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    128: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd127;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd150;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    129: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd128;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd128;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    130: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd130;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd68;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    131: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd131;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd150;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    132: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd132;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd132;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    133: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd133;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd68;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd68;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    134: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd136;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd8;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    135: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd134;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd150;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    136: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd138;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd156;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    137: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd68;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd68;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd68;
      21: stateTransition = 11'd136;
      22: stateTransition = 11'd68;
      23: stateTransition = 11'd68;
      24: stateTransition = 11'd68;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd68;
      27: stateTransition = 11'd68;
      28: stateTransition = 11'd68;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd68;
      31: stateTransition = 11'd68;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    138: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    139: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd154;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    140: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd142;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd148;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    141: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd143;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd148;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    142: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd144;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd148;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    143: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd145;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd148;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    144: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd146;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    145: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd148;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd148;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    146: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd148;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd148;
      19: stateTransition = 11'd148;
      20: stateTransition = 11'd148;
      21: stateTransition = 11'd146;
      22: stateTransition = 11'd148;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd148;
      25: stateTransition = 11'd148;
      26: stateTransition = 11'd148;
      27: stateTransition = 11'd148;
      28: stateTransition = 11'd148;
      29: stateTransition = 11'd148;
      30: stateTransition = 11'd148;
      31: stateTransition = 11'd148;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    147: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd150;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    148: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd138;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd150;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    149: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd141;
      2: stateTransition = 11'd141;
      3: stateTransition = 11'd141;
      4: stateTransition = 11'd147;
      5: stateTransition = 11'd141;
      6: stateTransition = 11'd93;
      7: stateTransition = 11'd141;
      8: stateTransition = 11'd141;
      9: stateTransition = 11'd141;
      10: stateTransition = 11'd141;
      11: stateTransition = 11'd141;
      12: stateTransition = 11'd141;
      13: stateTransition = 11'd141;
      14: stateTransition = 11'd141;
      15: stateTransition = 11'd141;
      16: stateTransition = 11'd141;
      17: stateTransition = 11'd141;
      18: stateTransition = 11'd141;
      19: stateTransition = 11'd141;
      20: stateTransition = 11'd141;
      21: stateTransition = 11'd141;
      22: stateTransition = 11'd141;
      23: stateTransition = 11'd141;
      24: stateTransition = 11'd141;
      25: stateTransition = 11'd141;
      26: stateTransition = 11'd141;
      27: stateTransition = 11'd141;
      28: stateTransition = 11'd141;
      29: stateTransition = 11'd141;
      30: stateTransition = 11'd141;
      31: stateTransition = 11'd141;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    150: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd150;
      19: stateTransition = 11'd150;
      20: stateTransition = 11'd150;
      21: stateTransition = 11'd150;
      22: stateTransition = 11'd150;
      23: stateTransition = 11'd150;
      24: stateTransition = 11'd156;
      25: stateTransition = 11'd150;
      26: stateTransition = 11'd150;
      27: stateTransition = 11'd150;
      28: stateTransition = 11'd150;
      29: stateTransition = 11'd150;
      30: stateTransition = 11'd150;
      31: stateTransition = 11'd150;
      32: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
