 count_ALL_0 ,
 count_ALL_1 ,
 count_ALL_2 ,
 count_ALL_3 ,
 count_ALL_4 ,
 count_finger_0 ,
 count_ftp_0 ,
 count_http_0 ,
 count_imap_0 ,
 count_netbios_0 ,
 count_nntp_0 ,
 count_pop3_0 ,
 count_rlogin_0 ,
 count_smtp_0 ,
 count_telnet_0 ,
 count_CATEGORY_finger ,
 count_CATEGORY_ftp ,
 count_CATEGORY_http ,
 count_CATEGORY_imap ,
 count_CATEGORY_netbios ,
 count_CATEGORY_nntp ,
 count_CATEGORY_pop3 ,
 count_CATEGORY_rlogin ,
 count_CATEGORY_smtp ,
 count_CATEGORY_telnet ,

`ifdef REGEX_OPTIONAL
count_ALL_5 ,
count_ALL_6 ,
count_ALL_7 ,
count_ALL_8 ,
count_ALL_9 ,
count_ALL_10 ,
count_ALL_11 ,
count_ALL_12 ,
count_ALL_13 ,
count_ALL_14 ,

count_finger_1 ,
count_finger_2 ,
count_finger_3 ,
count_finger_4 ,
count_finger_5 ,

count_ftp_1 ,
count_ftp_2 ,
count_ftp_3 ,
count_ftp_4 ,
count_ftp_5 ,
count_ftp_6 ,
count_ftp_7 ,
count_ftp_8 ,
count_ftp_9 ,



count_http_1 ,
count_http_2 ,
count_http_3 ,
count_http_4 ,
count_http_5 ,
count_http_6 ,
count_http_7 ,
count_http_8 ,
count_http_9 ,

count_imap_1 ,
count_imap_2 ,
count_imap_3 ,
count_imap_4 ,
count_imap_5 ,
count_imap_6 ,
count_imap_7 ,
count_imap_8 ,
count_imap_9 ,

count_netbios_1 ,
count_netbios_2 ,
count_netbios_3 ,
count_netbios_4 ,
count_netbios_5 ,
count_netbios_6 ,
count_netbios_7 ,
count_netbios_8 ,
count_netbios_9 ,

count_nntp_1 ,
count_nntp_2 ,
count_nntp_3 ,
count_nntp_4 ,
count_nntp_5 ,
count_nntp_6 ,
count_nntp_7 ,
count_nntp_8 ,
count_nntp_9 ,

count_pop3_1 ,
count_pop3_2 ,
count_pop3_3 ,
count_pop3_4 ,
count_pop3_5 ,
count_pop3_6 ,
count_pop3_7 ,
count_pop3_8 ,
count_pop3_9 ,


count_rlogin_1 ,
count_rlogin_2 ,
count_rlogin_3 ,
count_rlogin_4 ,
count_rlogin_5 ,


count_smtp_1 ,
count_smtp_2 ,
count_smtp_3 ,
count_smtp_4 ,
count_smtp_5 ,
count_smtp_6 ,
count_smtp_7 ,
count_smtp_8 ,
count_smtp_9 ,


count_telnet_1 ,
count_telnet_2 ,
count_telnet_3 ,
count_telnet_4 ,
count_telnet_5 ,
count_telnet_6 ,
count_telnet_7 ,
count_telnet_8 ,
count_telnet_9 ,

count_CATEGORY_aim ,
count_CATEGORY_bittorrent ,
count_CATEGORY_cvs ,
count_CATEGORY_dhcp ,
count_CATEGORY_directconnect ,
count_CATEGORY_dns ,
count_CATEGORY_fasttrack ,
count_CATEGORY_tor ,
count_CATEGORY_vnc ,
count_CATEGORY_worldofwarcraft ,
count_CATEGORY_x11 ,
count_CATEGORY_yahoo ,
count_CATEGORY_freenet ,
count_CATEGORY_gnutella ,
count_CATEGORY_gopher ,
count_CATEGORY_irc ,
count_CATEGORY_jabber ,
count_CATEGORY_msn ,
count_CATEGORY_napster ,
count_CATEGORY_sip ,
count_CATEGORY_snmp ,
count_CATEGORY_socks ,
count_CATEGORY_ssh ,
count_CATEGORY_ssl ,
count_CATEGORY_subversion ,    
`endif //  `ifdef REGEX_OPTIONAL
