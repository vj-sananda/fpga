`timescale 1ns/1ps

`define ENABLED_REGEX_http_6 TRUE

module http_6_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_http_6

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd16;
    1: charMap = 8'd16;
    2: charMap = 8'd16;
    3: charMap = 8'd16;
    4: charMap = 8'd16;
    5: charMap = 8'd16;
    6: charMap = 8'd16;
    7: charMap = 8'd16;
    8: charMap = 8'd16;
    9: charMap = 8'd11;
    10: charMap = 8'd12;
    11: charMap = 8'd11;
    12: charMap = 8'd16;
    13: charMap = 8'd11;
    14: charMap = 8'd16;
    15: charMap = 8'd16;
    16: charMap = 8'd16;
    17: charMap = 8'd16;
    18: charMap = 8'd16;
    19: charMap = 8'd16;
    20: charMap = 8'd16;
    21: charMap = 8'd16;
    22: charMap = 8'd16;
    23: charMap = 8'd16;
    24: charMap = 8'd16;
    25: charMap = 8'd16;
    26: charMap = 8'd16;
    27: charMap = 8'd16;
    28: charMap = 8'd16;
    29: charMap = 8'd16;
    30: charMap = 8'd16;
    31: charMap = 8'd16;
    32: charMap = 8'd11;
    33: charMap = 8'd16;
    34: charMap = 8'd16;
    35: charMap = 8'd16;
    36: charMap = 8'd16;
    37: charMap = 8'd16;
    38: charMap = 8'd16;
    39: charMap = 8'd16;
    40: charMap = 8'd16;
    41: charMap = 8'd16;
    42: charMap = 8'd16;
    43: charMap = 8'd16;
    44: charMap = 8'd16;
    45: charMap = 8'd16;
    46: charMap = 8'd16;
    47: charMap = 8'd16;
    48: charMap = 8'd16;
    49: charMap = 8'd16;
    50: charMap = 8'd16;
    51: charMap = 8'd16;
    52: charMap = 8'd16;
    53: charMap = 8'd16;
    54: charMap = 8'd16;
    55: charMap = 8'd16;
    56: charMap = 8'd16;
    57: charMap = 8'd16;
    58: charMap = 8'd10;
    59: charMap = 8'd16;
    60: charMap = 8'd16;
    61: charMap = 8'd16;
    62: charMap = 8'd16;
    63: charMap = 8'd16;
    64: charMap = 8'd16;
    65: charMap = 8'd1;
    66: charMap = 8'd13;
    67: charMap = 8'd15;
    68: charMap = 8'd16;
    69: charMap = 8'd16;
    70: charMap = 8'd16;
    71: charMap = 8'd16;
    72: charMap = 8'd4;
    73: charMap = 8'd7;
    74: charMap = 8'd16;
    75: charMap = 8'd16;
    76: charMap = 8'd16;
    77: charMap = 8'd16;
    78: charMap = 8'd9;
    79: charMap = 8'd5;
    80: charMap = 8'd16;
    81: charMap = 8'd16;
    82: charMap = 8'd6;
    83: charMap = 8'd14;
    84: charMap = 8'd3;
    85: charMap = 8'd2;
    86: charMap = 8'd16;
    87: charMap = 8'd16;
    88: charMap = 8'd16;
    89: charMap = 8'd16;
    90: charMap = 8'd8;
    91: charMap = 8'd16;
    92: charMap = 8'd16;
    93: charMap = 8'd16;
    94: charMap = 8'd16;
    95: charMap = 8'd16;
    96: charMap = 8'd16;
    97: charMap = 8'd1;
    98: charMap = 8'd13;
    99: charMap = 8'd15;
    100: charMap = 8'd16;
    101: charMap = 8'd16;
    102: charMap = 8'd16;
    103: charMap = 8'd16;
    104: charMap = 8'd4;
    105: charMap = 8'd7;
    106: charMap = 8'd16;
    107: charMap = 8'd16;
    108: charMap = 8'd16;
    109: charMap = 8'd16;
    110: charMap = 8'd9;
    111: charMap = 8'd5;
    112: charMap = 8'd16;
    113: charMap = 8'd16;
    114: charMap = 8'd6;
    115: charMap = 8'd14;
    116: charMap = 8'd3;
    117: charMap = 8'd2;
    118: charMap = 8'd16;
    119: charMap = 8'd16;
    120: charMap = 8'd16;
    121: charMap = 8'd16;
    122: charMap = 8'd8;
    123: charMap = 8'd16;
    124: charMap = 8'd16;
    125: charMap = 8'd16;
    126: charMap = 8'd16;
    127: charMap = 8'd16;
    128: charMap = 8'd16;
    129: charMap = 8'd16;
    130: charMap = 8'd16;
    131: charMap = 8'd16;
    132: charMap = 8'd16;
    133: charMap = 8'd16;
    134: charMap = 8'd16;
    135: charMap = 8'd16;
    136: charMap = 8'd16;
    137: charMap = 8'd16;
    138: charMap = 8'd16;
    139: charMap = 8'd16;
    140: charMap = 8'd16;
    141: charMap = 8'd16;
    142: charMap = 8'd16;
    143: charMap = 8'd16;
    144: charMap = 8'd16;
    145: charMap = 8'd16;
    146: charMap = 8'd16;
    147: charMap = 8'd16;
    148: charMap = 8'd16;
    149: charMap = 8'd16;
    150: charMap = 8'd16;
    151: charMap = 8'd16;
    152: charMap = 8'd16;
    153: charMap = 8'd16;
    154: charMap = 8'd16;
    155: charMap = 8'd16;
    156: charMap = 8'd16;
    157: charMap = 8'd16;
    158: charMap = 8'd16;
    159: charMap = 8'd16;
    160: charMap = 8'd16;
    161: charMap = 8'd16;
    162: charMap = 8'd16;
    163: charMap = 8'd16;
    164: charMap = 8'd16;
    165: charMap = 8'd16;
    166: charMap = 8'd16;
    167: charMap = 8'd16;
    168: charMap = 8'd16;
    169: charMap = 8'd16;
    170: charMap = 8'd16;
    171: charMap = 8'd16;
    172: charMap = 8'd16;
    173: charMap = 8'd16;
    174: charMap = 8'd16;
    175: charMap = 8'd16;
    176: charMap = 8'd16;
    177: charMap = 8'd16;
    178: charMap = 8'd16;
    179: charMap = 8'd16;
    180: charMap = 8'd16;
    181: charMap = 8'd16;
    182: charMap = 8'd16;
    183: charMap = 8'd16;
    184: charMap = 8'd16;
    185: charMap = 8'd16;
    186: charMap = 8'd16;
    187: charMap = 8'd16;
    188: charMap = 8'd16;
    189: charMap = 8'd16;
    190: charMap = 8'd16;
    191: charMap = 8'd16;
    192: charMap = 8'd16;
    193: charMap = 8'd16;
    194: charMap = 8'd16;
    195: charMap = 8'd16;
    196: charMap = 8'd16;
    197: charMap = 8'd16;
    198: charMap = 8'd16;
    199: charMap = 8'd16;
    200: charMap = 8'd16;
    201: charMap = 8'd16;
    202: charMap = 8'd16;
    203: charMap = 8'd16;
    204: charMap = 8'd16;
    205: charMap = 8'd16;
    206: charMap = 8'd16;
    207: charMap = 8'd16;
    208: charMap = 8'd16;
    209: charMap = 8'd16;
    210: charMap = 8'd16;
    211: charMap = 8'd16;
    212: charMap = 8'd16;
    213: charMap = 8'd16;
    214: charMap = 8'd16;
    215: charMap = 8'd16;
    216: charMap = 8'd16;
    217: charMap = 8'd16;
    218: charMap = 8'd16;
    219: charMap = 8'd16;
    220: charMap = 8'd16;
    221: charMap = 8'd16;
    222: charMap = 8'd16;
    223: charMap = 8'd16;
    224: charMap = 8'd16;
    225: charMap = 8'd16;
    226: charMap = 8'd16;
    227: charMap = 8'd16;
    228: charMap = 8'd16;
    229: charMap = 8'd16;
    230: charMap = 8'd16;
    231: charMap = 8'd16;
    232: charMap = 8'd16;
    233: charMap = 8'd16;
    234: charMap = 8'd16;
    235: charMap = 8'd16;
    236: charMap = 8'd16;
    237: charMap = 8'd16;
    238: charMap = 8'd16;
    239: charMap = 8'd16;
    240: charMap = 8'd16;
    241: charMap = 8'd16;
    242: charMap = 8'd16;
    243: charMap = 8'd16;
    244: charMap = 8'd16;
    245: charMap = 8'd16;
    246: charMap = 8'd16;
    247: charMap = 8'd16;
    248: charMap = 8'd16;
    249: charMap = 8'd16;
    250: charMap = 8'd16;
    251: charMap = 8'd16;
    252: charMap = 8'd16;
    253: charMap = 8'd16;
    254: charMap = 8'd16;
    255: charMap = 8'd16;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd1;
    3: stateMap = 11'd2;
    4: stateMap = 11'd3;
    5: stateMap = 11'd4;
    6: stateMap = 11'd5;
    7: stateMap = 11'd6;
    8: stateMap = 11'd7;
    9: stateMap = 11'd8;
    10: stateMap = 11'd9;
    11: stateMap = 11'd10;
    12: stateMap = 11'd11;
    13: stateMap = 11'd12;
    14: stateMap = 11'd13;
    15: stateMap = 11'd14;
    16: stateMap = 11'd15;
    17: stateMap = 11'd16;
    18: stateMap = 11'd17;
    19: stateMap = 11'd18;
    20: stateMap = 11'd19;
    21: stateMap = 11'd20;
    22: stateMap = 11'd21;
    23: stateMap = 11'd22;
    24: stateMap = 11'd23;
    25: stateMap = 11'd24;
    26: stateMap = 11'd25;
    27: stateMap = 11'd26;
    28: stateMap = 11'd27;
    29: stateMap = 11'd28;
    30: stateMap = 11'd29;
    31: stateMap = 11'd30;
    32: stateMap = 11'd31;
    33: stateMap = 11'd32;
    34: stateMap = 11'd33;
    35: stateMap = 11'd34;
    36: stateMap = 11'd35;
    37: stateMap = 11'd36;
    38: stateMap = 11'd37;
    39: stateMap = 11'd38;
    40: stateMap = 11'd39;
    41: stateMap = 11'd40;
    42: stateMap = 11'd41;
    43: stateMap = 11'd42;
    44: stateMap = 11'd43;
    45: stateMap = 11'd44;
    46: stateMap = 11'd45;
    47: stateMap = 11'd46;
    48: stateMap = 11'd47;
    49: stateMap = 11'd48;
    50: stateMap = 11'd49;
    51: stateMap = 11'd50;
    52: stateMap = 11'd51;
    53: stateMap = 11'd52;
    54: stateMap = 11'd53;
    55: stateMap = 11'd54;
    56: stateMap = 11'd55;
    57: stateMap = 11'd56;
    58: stateMap = 11'd57;
    59: stateMap = 11'd58;
    60: stateMap = 11'd59;
    61: stateMap = 11'd60;
    62: stateMap = 11'd61;
    63: stateMap = 11'd62;
    64: stateMap = 11'd63;
    65: stateMap = 11'd64;
    66: stateMap = 11'd65;
    67: stateMap = 11'd66;
    68: stateMap = 11'd67;
    69: stateMap = 11'd68;
    70: stateMap = 11'd69;
    71: stateMap = 11'd70;
    72: stateMap = 11'd71;
    73: stateMap = 11'd72;
    74: stateMap = 11'd73;
    75: stateMap = 11'd74;
    76: stateMap = 11'd75;
    77: stateMap = 11'd76;
    78: stateMap = 11'd77;
    79: stateMap = 11'd78;
    80: stateMap = 11'd79;
    81: stateMap = 11'd80;
    82: stateMap = 11'd81;
    83: stateMap = 11'd82;
    84: stateMap = 11'd83;
    85: stateMap = 11'd84;
    86: stateMap = 11'd85;
    87: stateMap = 11'd86;
    88: stateMap = 11'd87;
    89: stateMap = 11'd88;
    90: stateMap = 11'd89;
    91: stateMap = 11'd90;
    92: stateMap = 11'd91;
    93: stateMap = 11'd92;
    94: stateMap = 11'd93;
    95: stateMap = 11'd94;
    96: stateMap = 11'd95;
    97: stateMap = 11'd96;
    98: stateMap = 11'd97;
    99: stateMap = 11'd98;
    100: stateMap = 11'd99;
    101: stateMap = 11'd100;
    102: stateMap = 11'd101;
    103: stateMap = 11'd102;
    104: stateMap = 11'd103;
    105: stateMap = 11'd104;
    106: stateMap = 11'd105;
    107: stateMap = 11'd106;
    108: stateMap = 11'd107;
    109: stateMap = 11'd108;
    110: stateMap = 11'd109;
    111: stateMap = 11'd110;
    112: stateMap = 11'd111;
    113: stateMap = 11'd112;
    114: stateMap = 11'd113;
    115: stateMap = 11'd114;
    116: stateMap = 11'd115;
    117: stateMap = 11'd116;
    118: stateMap = 11'd117;
    119: stateMap = 11'd118;
    120: stateMap = 11'd119;
    121: stateMap = 11'd120;
    122: stateMap = 11'd121;
    123: stateMap = 11'd122;
    124: stateMap = 11'd123;
    125: stateMap = 11'd124;
    126: stateMap = 11'd125;
    127: stateMap = 11'd126;
    128: stateMap = 11'd127;
    129: stateMap = 11'd128;
    130: stateMap = 11'd129;
    131: stateMap = 11'd130;
    132: stateMap = 11'd131;
    133: stateMap = 11'd132;
    134: stateMap = 11'd133;
    135: stateMap = 11'd134;
    136: stateMap = 11'd135;
    137: stateMap = 11'd136;
    138: stateMap = 11'd137;
    139: stateMap = 11'd138;
    140: stateMap = 11'd139;
    141: stateMap = 11'd140;
    142: stateMap = 11'd141;
    143: stateMap = 11'd142;
    144: stateMap = 11'd143;
    145: stateMap = 11'd144;
    146: stateMap = 11'd145;
    147: stateMap = 11'd146;
    148: stateMap = 11'd147;
    149: stateMap = 11'd148;
    150: stateMap = 11'd149;
    151: stateMap = 11'd150;
    152: stateMap = 11'd151;
    153: stateMap = 11'd152;
    154: stateMap = 11'd153;
    155: stateMap = 11'd154;
    156: stateMap = 11'd155;
    157: stateMap = 11'd156;
    158: stateMap = 11'd157;
    159: stateMap = 11'd158;
    160: stateMap = 11'd159;
    161: stateMap = 11'd160;
    162: stateMap = 11'd161;
    163: stateMap = 11'd162;
    164: stateMap = 11'd163;
    165: stateMap = 11'd164;
    166: stateMap = 11'd165;
    167: stateMap = 11'd166;
    168: stateMap = 11'd167;
    169: stateMap = 11'd168;
    170: stateMap = 11'd169;
    171: stateMap = 11'd170;
    172: stateMap = 11'd171;
    173: stateMap = 11'd172;
    174: stateMap = 11'd173;
    175: stateMap = 11'd174;
    176: stateMap = 11'd175;
    177: stateMap = 11'd176;
    178: stateMap = 11'd177;
    179: stateMap = 11'd178;
    180: stateMap = 11'd179;
    181: stateMap = 11'd180;
    182: stateMap = 11'd181;
    183: stateMap = 11'd182;
    184: stateMap = 11'd183;
    185: stateMap = 11'd184;
    186: stateMap = 11'd185;
    187: stateMap = 11'd186;
    188: stateMap = 11'd187;
    189: stateMap = 11'd188;
    190: stateMap = 11'd189;
    191: stateMap = 11'd190;
    192: stateMap = 11'd191;
    193: stateMap = 11'd192;
    194: stateMap = 11'd193;
    195: stateMap = 11'd194;
    196: stateMap = 11'd195;
    197: stateMap = 11'd196;
    198: stateMap = 11'd197;
    199: stateMap = 11'd198;
    200: stateMap = 11'd199;
    201: stateMap = 11'd200;
    202: stateMap = 11'd201;
    203: stateMap = 11'd202;
    204: stateMap = 11'd203;
    205: stateMap = 11'd204;
    206: stateMap = 11'd205;
    207: stateMap = 11'd206;
    208: stateMap = 11'd207;
    209: stateMap = 11'd208;
    210: stateMap = 11'd209;
    211: stateMap = 11'd210;
    212: stateMap = 11'd211;
    213: stateMap = 11'd212;
    214: stateMap = 11'd213;
    215: stateMap = 11'd214;
    216: stateMap = 11'd215;
    217: stateMap = 11'd216;
    218: stateMap = 11'd217;
    219: stateMap = 11'd218;
    220: stateMap = 11'd219;
    221: stateMap = 11'd220;
    222: stateMap = 11'd221;
    223: stateMap = 11'd222;
    224: stateMap = 11'd223;
    225: stateMap = 11'd224;
    226: stateMap = 11'd225;
    227: stateMap = 11'd226;
    228: stateMap = 11'd227;
    229: stateMap = 11'd228;
    230: stateMap = 11'd229;
    231: stateMap = 11'd230;
    232: stateMap = 11'd231;
    233: stateMap = 11'd232;
    234: stateMap = 11'd233;
    235: stateMap = 11'd234;
    236: stateMap = 11'd235;
    237: stateMap = 11'd236;
    238: stateMap = 11'd237;
    239: stateMap = 11'd238;
    240: stateMap = 11'd239;
    241: stateMap = 11'd240;
    242: stateMap = 11'd241;
    243: stateMap = 11'd242;
    244: stateMap = 11'd243;
    245: stateMap = 11'd244;
    246: stateMap = 11'd245;
    247: stateMap = 11'd246;
    248: stateMap = 11'd247;
    249: stateMap = 11'd248;
    250: stateMap = 11'd249;
    251: stateMap = 11'd250;
    252: stateMap = 11'd251;
    253: stateMap = 11'd252;
    254: stateMap = 11'd253;
    255: stateMap = 11'd254;
    256: stateMap = 11'd255;
    257: stateMap = 11'd256;
    258: stateMap = 11'd257;
    259: stateMap = 11'd258;
    260: stateMap = 11'd259;
    261: stateMap = 11'd260;
    262: stateMap = 11'd261;
    263: stateMap = 11'd262;
    264: stateMap = 11'd263;
    265: stateMap = 11'd264;
    266: stateMap = 11'd265;
    267: stateMap = 11'd266;
    268: stateMap = 11'd267;
    269: stateMap = 11'd268;
    270: stateMap = 11'd269;
    271: stateMap = 11'd270;
    272: stateMap = 11'd271;
    273: stateMap = 11'd272;
    274: stateMap = 11'd273;
    275: stateMap = 11'd274;
    276: stateMap = 11'd275;
    277: stateMap = 11'd276;
    278: stateMap = 11'd277;
    279: stateMap = 11'd278;
    280: stateMap = 11'd279;
    281: stateMap = 11'd280;
    282: stateMap = 11'd281;
    283: stateMap = 11'd282;
    284: stateMap = 11'd283;
    285: stateMap = 11'd284;
    286: stateMap = 11'd285;
    287: stateMap = 11'd286;
    288: stateMap = 11'd287;
    289: stateMap = 11'd288;
    290: stateMap = 11'd289;
    291: stateMap = 11'd290;
    292: stateMap = 11'd291;
    293: stateMap = 11'd292;
    294: stateMap = 11'd293;
    295: stateMap = 11'd294;
    296: stateMap = 11'd295;
    297: stateMap = 11'd296;
    298: stateMap = 11'd297;
    299: stateMap = 11'd298;
    300: stateMap = 11'd299;
    301: stateMap = 11'd300;
    302: stateMap = 11'd301;
    303: stateMap = 11'd302;
    304: stateMap = 11'd303;
    305: stateMap = 11'd304;
    306: stateMap = 11'd305;
    307: stateMap = 11'd306;
    308: stateMap = 11'd307;
    309: stateMap = 11'd308;
    310: stateMap = 11'd309;
    311: stateMap = 11'd310;
    312: stateMap = 11'd311;
    313: stateMap = 11'd312;
    314: stateMap = 11'd313;
    315: stateMap = 11'd314;
    316: stateMap = 11'd315;
    317: stateMap = 11'd316;
    318: stateMap = 11'd317;
    319: stateMap = 11'd318;
    320: stateMap = 11'd319;
    321: stateMap = 11'd320;
    322: stateMap = 11'd321;
    323: stateMap = 11'd322;
    324: stateMap = 11'd323;
    325: stateMap = 11'd324;
    326: stateMap = 11'd325;
    327: stateMap = 11'd326;
    328: stateMap = 11'd327;
    329: stateMap = 11'd328;
    330: stateMap = 11'd329;
    331: stateMap = 11'd330;
    332: stateMap = 11'd331;
    333: stateMap = 11'd332;
    334: stateMap = 11'd333;
    335: stateMap = 11'd334;
    336: stateMap = 11'd335;
    337: stateMap = 11'd336;
    338: stateMap = 11'd337;
    339: stateMap = 11'd338;
    340: stateMap = 11'd339;
    341: stateMap = 11'd340;
    342: stateMap = 11'd341;
    343: stateMap = 11'd342;
    344: stateMap = 11'd343;
    345: stateMap = 11'd344;
    346: stateMap = 11'd345;
    347: stateMap = 11'd346;
    348: stateMap = 11'd347;
    349: stateMap = 11'd348;
    350: stateMap = 11'd349;
    351: stateMap = 11'd350;
    352: stateMap = 11'd351;
    353: stateMap = 11'd352;
    354: stateMap = 11'd353;
    355: stateMap = 11'd354;
    356: stateMap = 11'd355;
    357: stateMap = 11'd356;
    358: stateMap = 11'd357;
    359: stateMap = 11'd358;
    360: stateMap = 11'd359;
    361: stateMap = 11'd360;
    362: stateMap = 11'd361;
    363: stateMap = 11'd362;
    364: stateMap = 11'd363;
    365: stateMap = 11'd364;
    366: stateMap = 11'd365;
    367: stateMap = 11'd366;
    368: stateMap = 11'd367;
    369: stateMap = 11'd368;
    370: stateMap = 11'd369;
    371: stateMap = 11'd370;
    372: stateMap = 11'd371;
    373: stateMap = 11'd372;
    374: stateMap = 11'd373;
    375: stateMap = 11'd374;
    376: stateMap = 11'd375;
    377: stateMap = 11'd376;
    378: stateMap = 11'd377;
    379: stateMap = 11'd378;
    380: stateMap = 11'd379;
    381: stateMap = 11'd380;
    382: stateMap = 11'd381;
    383: stateMap = 11'd382;
    384: stateMap = 11'd383;
    385: stateMap = 11'd384;
    386: stateMap = 11'd385;
    387: stateMap = 11'd386;
    388: stateMap = 11'd387;
    389: stateMap = 11'd388;
    390: stateMap = 11'd389;
    391: stateMap = 11'd390;
    392: stateMap = 11'd391;
    393: stateMap = 11'd392;
    394: stateMap = 11'd393;
    395: stateMap = 11'd394;
    396: stateMap = 11'd395;
    397: stateMap = 11'd396;
    398: stateMap = 11'd397;
    399: stateMap = 11'd398;
    400: stateMap = 11'd399;
    401: stateMap = 11'd400;
    402: stateMap = 11'd401;
    403: stateMap = 11'd402;
    404: stateMap = 11'd403;
    405: stateMap = 11'd404;
    406: stateMap = 11'd405;
    407: stateMap = 11'd406;
    408: stateMap = 11'd407;
    409: stateMap = 11'd408;
    410: stateMap = 11'd409;
    411: stateMap = 11'd410;
    412: stateMap = 11'd411;
    413: stateMap = 11'd412;
    414: stateMap = 11'd413;
    415: stateMap = 11'd414;
    416: stateMap = 11'd415;
    417: stateMap = 11'd416;
    418: stateMap = 11'd417;
    419: stateMap = 11'd418;
    420: stateMap = 11'd419;
    421: stateMap = 11'd420;
    422: stateMap = 11'd421;
    423: stateMap = 11'd422;
    424: stateMap = 11'd423;
    425: stateMap = 11'd424;
    426: stateMap = 11'd425;
    427: stateMap = 11'd426;
    428: stateMap = 11'd427;
    429: stateMap = 11'd428;
    430: stateMap = 11'd429;
    431: stateMap = 11'd430;
    432: stateMap = 11'd431;
    433: stateMap = 11'd432;
    434: stateMap = 11'd433;
    435: stateMap = 11'd434;
    436: stateMap = 11'd435;
    437: stateMap = 11'd436;
    438: stateMap = 11'd437;
    439: stateMap = 11'd438;
    440: stateMap = 11'd439;
    441: stateMap = 11'd440;
    442: stateMap = 11'd441;
    443: stateMap = 11'd442;
    444: stateMap = 11'd443;
    445: stateMap = 11'd444;
    446: stateMap = 11'd445;
    447: stateMap = 11'd446;
    448: stateMap = 11'd447;
    449: stateMap = 11'd448;
    450: stateMap = 11'd449;
    451: stateMap = 11'd450;
    452: stateMap = 11'd451;
    453: stateMap = 11'd452;
    454: stateMap = 11'd453;
    455: stateMap = 11'd454;
    456: stateMap = 11'd455;
    457: stateMap = 11'd456;
    458: stateMap = 11'd457;
    459: stateMap = 11'd458;
    460: stateMap = 11'd459;
    461: stateMap = 11'd460;
    462: stateMap = 11'd461;
    463: stateMap = 11'd462;
    464: stateMap = 11'd463;
    465: stateMap = 11'd464;
    466: stateMap = 11'd465;
    467: stateMap = 11'd466;
    468: stateMap = 11'd467;
    469: stateMap = 11'd468;
    470: stateMap = 11'd469;
    471: stateMap = 11'd470;
    472: stateMap = 11'd471;
    473: stateMap = 11'd472;
    474: stateMap = 11'd473;
    475: stateMap = 11'd474;
    476: stateMap = 11'd475;
    477: stateMap = 11'd476;
    478: stateMap = 11'd477;
    479: stateMap = 11'd478;
    480: stateMap = 11'd479;
    481: stateMap = 11'd480;
    482: stateMap = 11'd481;
    483: stateMap = 11'd482;
    484: stateMap = 11'd483;
    485: stateMap = 11'd484;
    486: stateMap = 11'd485;
    487: stateMap = 11'd486;
    488: stateMap = 11'd487;
    489: stateMap = 11'd488;
    490: stateMap = 11'd489;
    491: stateMap = 11'd490;
    492: stateMap = 11'd491;
    493: stateMap = 11'd492;
    494: stateMap = 11'd493;
    495: stateMap = 11'd494;
    496: stateMap = 11'd495;
    497: stateMap = 11'd496;
    498: stateMap = 11'd497;
    499: stateMap = 11'd498;
    500: stateMap = 11'd499;
    501: stateMap = 11'd500;
    502: stateMap = 11'd501;
    503: stateMap = 11'd502;
    504: stateMap = 11'd503;
    505: stateMap = 11'd504;
    506: stateMap = 11'd505;
    507: stateMap = 11'd506;
    508: stateMap = 11'd507;
    509: stateMap = 11'd508;
    510: stateMap = 11'd509;
    511: stateMap = 11'd510;
    512: stateMap = 11'd511;
    513: stateMap = 11'd512;
    514: stateMap = 11'd513;
    515: stateMap = 11'd514;
    516: stateMap = 11'd515;
    517: stateMap = 11'd516;
    518: stateMap = 11'd517;
    519: stateMap = 11'd518;
    520: stateMap = 11'd519;
    521: stateMap = 11'd520;
    522: stateMap = 11'd521;
    523: stateMap = 11'd522;
    524: stateMap = 11'd523;
    525: stateMap = 11'd524;
    526: stateMap = 11'd525;
    527: stateMap = 11'd526;
    528: stateMap = 11'd527;
    529: stateMap = 11'd528;
    530: stateMap = 11'd529;
    531: stateMap = 11'd530;
    532: stateMap = 11'd531;
    533: stateMap = 11'd532;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b0;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b0;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b0;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b0;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b0;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b0;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b0;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b0;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b0;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b0;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b0;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b0;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b0;
    62: acceptStates = 1'b0;
    63: acceptStates = 1'b0;
    64: acceptStates = 1'b0;
    65: acceptStates = 1'b0;
    66: acceptStates = 1'b0;
    67: acceptStates = 1'b0;
    68: acceptStates = 1'b0;
    69: acceptStates = 1'b0;
    70: acceptStates = 1'b0;
    71: acceptStates = 1'b0;
    72: acceptStates = 1'b0;
    73: acceptStates = 1'b0;
    74: acceptStates = 1'b0;
    75: acceptStates = 1'b0;
    76: acceptStates = 1'b0;
    77: acceptStates = 1'b0;
    78: acceptStates = 1'b0;
    79: acceptStates = 1'b0;
    80: acceptStates = 1'b0;
    81: acceptStates = 1'b0;
    82: acceptStates = 1'b0;
    83: acceptStates = 1'b0;
    84: acceptStates = 1'b0;
    85: acceptStates = 1'b0;
    86: acceptStates = 1'b0;
    87: acceptStates = 1'b0;
    88: acceptStates = 1'b0;
    89: acceptStates = 1'b0;
    90: acceptStates = 1'b0;
    91: acceptStates = 1'b0;
    92: acceptStates = 1'b0;
    93: acceptStates = 1'b0;
    94: acceptStates = 1'b0;
    95: acceptStates = 1'b0;
    96: acceptStates = 1'b0;
    97: acceptStates = 1'b0;
    98: acceptStates = 1'b0;
    99: acceptStates = 1'b0;
    100: acceptStates = 1'b0;
    101: acceptStates = 1'b0;
    102: acceptStates = 1'b0;
    103: acceptStates = 1'b0;
    104: acceptStates = 1'b0;
    105: acceptStates = 1'b0;
    106: acceptStates = 1'b0;
    107: acceptStates = 1'b0;
    108: acceptStates = 1'b0;
    109: acceptStates = 1'b0;
    110: acceptStates = 1'b0;
    111: acceptStates = 1'b0;
    112: acceptStates = 1'b0;
    113: acceptStates = 1'b0;
    114: acceptStates = 1'b0;
    115: acceptStates = 1'b0;
    116: acceptStates = 1'b0;
    117: acceptStates = 1'b0;
    118: acceptStates = 1'b0;
    119: acceptStates = 1'b0;
    120: acceptStates = 1'b0;
    121: acceptStates = 1'b0;
    122: acceptStates = 1'b0;
    123: acceptStates = 1'b0;
    124: acceptStates = 1'b0;
    125: acceptStates = 1'b0;
    126: acceptStates = 1'b0;
    127: acceptStates = 1'b0;
    128: acceptStates = 1'b0;
    129: acceptStates = 1'b0;
    130: acceptStates = 1'b0;
    131: acceptStates = 1'b0;
    132: acceptStates = 1'b0;
    133: acceptStates = 1'b0;
    134: acceptStates = 1'b0;
    135: acceptStates = 1'b0;
    136: acceptStates = 1'b0;
    137: acceptStates = 1'b0;
    138: acceptStates = 1'b0;
    139: acceptStates = 1'b0;
    140: acceptStates = 1'b0;
    141: acceptStates = 1'b0;
    142: acceptStates = 1'b0;
    143: acceptStates = 1'b0;
    144: acceptStates = 1'b0;
    145: acceptStates = 1'b0;
    146: acceptStates = 1'b0;
    147: acceptStates = 1'b0;
    148: acceptStates = 1'b0;
    149: acceptStates = 1'b0;
    150: acceptStates = 1'b0;
    151: acceptStates = 1'b0;
    152: acceptStates = 1'b0;
    153: acceptStates = 1'b0;
    154: acceptStates = 1'b0;
    155: acceptStates = 1'b0;
    156: acceptStates = 1'b0;
    157: acceptStates = 1'b0;
    158: acceptStates = 1'b0;
    159: acceptStates = 1'b0;
    160: acceptStates = 1'b0;
    161: acceptStates = 1'b0;
    162: acceptStates = 1'b0;
    163: acceptStates = 1'b0;
    164: acceptStates = 1'b0;
    165: acceptStates = 1'b0;
    166: acceptStates = 1'b0;
    167: acceptStates = 1'b0;
    168: acceptStates = 1'b0;
    169: acceptStates = 1'b0;
    170: acceptStates = 1'b0;
    171: acceptStates = 1'b0;
    172: acceptStates = 1'b0;
    173: acceptStates = 1'b0;
    174: acceptStates = 1'b0;
    175: acceptStates = 1'b0;
    176: acceptStates = 1'b0;
    177: acceptStates = 1'b0;
    178: acceptStates = 1'b0;
    179: acceptStates = 1'b0;
    180: acceptStates = 1'b0;
    181: acceptStates = 1'b0;
    182: acceptStates = 1'b0;
    183: acceptStates = 1'b0;
    184: acceptStates = 1'b0;
    185: acceptStates = 1'b0;
    186: acceptStates = 1'b0;
    187: acceptStates = 1'b0;
    188: acceptStates = 1'b0;
    189: acceptStates = 1'b0;
    190: acceptStates = 1'b0;
    191: acceptStates = 1'b0;
    192: acceptStates = 1'b0;
    193: acceptStates = 1'b0;
    194: acceptStates = 1'b0;
    195: acceptStates = 1'b0;
    196: acceptStates = 1'b0;
    197: acceptStates = 1'b0;
    198: acceptStates = 1'b0;
    199: acceptStates = 1'b0;
    200: acceptStates = 1'b0;
    201: acceptStates = 1'b0;
    202: acceptStates = 1'b0;
    203: acceptStates = 1'b0;
    204: acceptStates = 1'b0;
    205: acceptStates = 1'b0;
    206: acceptStates = 1'b0;
    207: acceptStates = 1'b0;
    208: acceptStates = 1'b0;
    209: acceptStates = 1'b0;
    210: acceptStates = 1'b0;
    211: acceptStates = 1'b0;
    212: acceptStates = 1'b0;
    213: acceptStates = 1'b0;
    214: acceptStates = 1'b0;
    215: acceptStates = 1'b0;
    216: acceptStates = 1'b0;
    217: acceptStates = 1'b0;
    218: acceptStates = 1'b0;
    219: acceptStates = 1'b0;
    220: acceptStates = 1'b0;
    221: acceptStates = 1'b0;
    222: acceptStates = 1'b0;
    223: acceptStates = 1'b0;
    224: acceptStates = 1'b0;
    225: acceptStates = 1'b0;
    226: acceptStates = 1'b0;
    227: acceptStates = 1'b0;
    228: acceptStates = 1'b0;
    229: acceptStates = 1'b0;
    230: acceptStates = 1'b0;
    231: acceptStates = 1'b0;
    232: acceptStates = 1'b0;
    233: acceptStates = 1'b0;
    234: acceptStates = 1'b0;
    235: acceptStates = 1'b0;
    236: acceptStates = 1'b0;
    237: acceptStates = 1'b0;
    238: acceptStates = 1'b0;
    239: acceptStates = 1'b0;
    240: acceptStates = 1'b0;
    241: acceptStates = 1'b0;
    242: acceptStates = 1'b0;
    243: acceptStates = 1'b0;
    244: acceptStates = 1'b0;
    245: acceptStates = 1'b0;
    246: acceptStates = 1'b0;
    247: acceptStates = 1'b0;
    248: acceptStates = 1'b0;
    249: acceptStates = 1'b0;
    250: acceptStates = 1'b0;
    251: acceptStates = 1'b0;
    252: acceptStates = 1'b0;
    253: acceptStates = 1'b0;
    254: acceptStates = 1'b0;
    255: acceptStates = 1'b0;
    256: acceptStates = 1'b0;
    257: acceptStates = 1'b0;
    258: acceptStates = 1'b0;
    259: acceptStates = 1'b0;
    260: acceptStates = 1'b0;
    261: acceptStates = 1'b0;
    262: acceptStates = 1'b0;
    263: acceptStates = 1'b0;
    264: acceptStates = 1'b0;
    265: acceptStates = 1'b0;
    266: acceptStates = 1'b0;
    267: acceptStates = 1'b0;
    268: acceptStates = 1'b0;
    269: acceptStates = 1'b0;
    270: acceptStates = 1'b0;
    271: acceptStates = 1'b0;
    272: acceptStates = 1'b0;
    273: acceptStates = 1'b0;
    274: acceptStates = 1'b0;
    275: acceptStates = 1'b0;
    276: acceptStates = 1'b0;
    277: acceptStates = 1'b0;
    278: acceptStates = 1'b0;
    279: acceptStates = 1'b0;
    280: acceptStates = 1'b0;
    281: acceptStates = 1'b0;
    282: acceptStates = 1'b0;
    283: acceptStates = 1'b0;
    284: acceptStates = 1'b0;
    285: acceptStates = 1'b0;
    286: acceptStates = 1'b0;
    287: acceptStates = 1'b0;
    288: acceptStates = 1'b0;
    289: acceptStates = 1'b0;
    290: acceptStates = 1'b0;
    291: acceptStates = 1'b0;
    292: acceptStates = 1'b0;
    293: acceptStates = 1'b0;
    294: acceptStates = 1'b0;
    295: acceptStates = 1'b0;
    296: acceptStates = 1'b0;
    297: acceptStates = 1'b0;
    298: acceptStates = 1'b0;
    299: acceptStates = 1'b0;
    300: acceptStates = 1'b0;
    301: acceptStates = 1'b0;
    302: acceptStates = 1'b0;
    303: acceptStates = 1'b0;
    304: acceptStates = 1'b0;
    305: acceptStates = 1'b0;
    306: acceptStates = 1'b0;
    307: acceptStates = 1'b0;
    308: acceptStates = 1'b0;
    309: acceptStates = 1'b0;
    310: acceptStates = 1'b0;
    311: acceptStates = 1'b0;
    312: acceptStates = 1'b0;
    313: acceptStates = 1'b0;
    314: acceptStates = 1'b0;
    315: acceptStates = 1'b0;
    316: acceptStates = 1'b0;
    317: acceptStates = 1'b0;
    318: acceptStates = 1'b0;
    319: acceptStates = 1'b0;
    320: acceptStates = 1'b0;
    321: acceptStates = 1'b0;
    322: acceptStates = 1'b0;
    323: acceptStates = 1'b0;
    324: acceptStates = 1'b0;
    325: acceptStates = 1'b0;
    326: acceptStates = 1'b0;
    327: acceptStates = 1'b0;
    328: acceptStates = 1'b0;
    329: acceptStates = 1'b0;
    330: acceptStates = 1'b0;
    331: acceptStates = 1'b0;
    332: acceptStates = 1'b0;
    333: acceptStates = 1'b0;
    334: acceptStates = 1'b0;
    335: acceptStates = 1'b0;
    336: acceptStates = 1'b0;
    337: acceptStates = 1'b0;
    338: acceptStates = 1'b0;
    339: acceptStates = 1'b0;
    340: acceptStates = 1'b0;
    341: acceptStates = 1'b0;
    342: acceptStates = 1'b0;
    343: acceptStates = 1'b0;
    344: acceptStates = 1'b0;
    345: acceptStates = 1'b0;
    346: acceptStates = 1'b0;
    347: acceptStates = 1'b0;
    348: acceptStates = 1'b0;
    349: acceptStates = 1'b0;
    350: acceptStates = 1'b0;
    351: acceptStates = 1'b0;
    352: acceptStates = 1'b0;
    353: acceptStates = 1'b0;
    354: acceptStates = 1'b0;
    355: acceptStates = 1'b0;
    356: acceptStates = 1'b0;
    357: acceptStates = 1'b0;
    358: acceptStates = 1'b0;
    359: acceptStates = 1'b0;
    360: acceptStates = 1'b0;
    361: acceptStates = 1'b0;
    362: acceptStates = 1'b0;
    363: acceptStates = 1'b0;
    364: acceptStates = 1'b0;
    365: acceptStates = 1'b0;
    366: acceptStates = 1'b0;
    367: acceptStates = 1'b0;
    368: acceptStates = 1'b0;
    369: acceptStates = 1'b0;
    370: acceptStates = 1'b0;
    371: acceptStates = 1'b0;
    372: acceptStates = 1'b0;
    373: acceptStates = 1'b0;
    374: acceptStates = 1'b0;
    375: acceptStates = 1'b0;
    376: acceptStates = 1'b0;
    377: acceptStates = 1'b0;
    378: acceptStates = 1'b0;
    379: acceptStates = 1'b0;
    380: acceptStates = 1'b0;
    381: acceptStates = 1'b0;
    382: acceptStates = 1'b0;
    383: acceptStates = 1'b0;
    384: acceptStates = 1'b0;
    385: acceptStates = 1'b0;
    386: acceptStates = 1'b0;
    387: acceptStates = 1'b0;
    388: acceptStates = 1'b0;
    389: acceptStates = 1'b0;
    390: acceptStates = 1'b0;
    391: acceptStates = 1'b0;
    392: acceptStates = 1'b0;
    393: acceptStates = 1'b0;
    394: acceptStates = 1'b0;
    395: acceptStates = 1'b0;
    396: acceptStates = 1'b0;
    397: acceptStates = 1'b0;
    398: acceptStates = 1'b0;
    399: acceptStates = 1'b0;
    400: acceptStates = 1'b0;
    401: acceptStates = 1'b0;
    402: acceptStates = 1'b0;
    403: acceptStates = 1'b0;
    404: acceptStates = 1'b0;
    405: acceptStates = 1'b0;
    406: acceptStates = 1'b0;
    407: acceptStates = 1'b0;
    408: acceptStates = 1'b0;
    409: acceptStates = 1'b0;
    410: acceptStates = 1'b0;
    411: acceptStates = 1'b0;
    412: acceptStates = 1'b0;
    413: acceptStates = 1'b0;
    414: acceptStates = 1'b0;
    415: acceptStates = 1'b0;
    416: acceptStates = 1'b0;
    417: acceptStates = 1'b0;
    418: acceptStates = 1'b0;
    419: acceptStates = 1'b0;
    420: acceptStates = 1'b0;
    421: acceptStates = 1'b0;
    422: acceptStates = 1'b0;
    423: acceptStates = 1'b0;
    424: acceptStates = 1'b0;
    425: acceptStates = 1'b0;
    426: acceptStates = 1'b0;
    427: acceptStates = 1'b0;
    428: acceptStates = 1'b0;
    429: acceptStates = 1'b0;
    430: acceptStates = 1'b0;
    431: acceptStates = 1'b0;
    432: acceptStates = 1'b0;
    433: acceptStates = 1'b0;
    434: acceptStates = 1'b0;
    435: acceptStates = 1'b0;
    436: acceptStates = 1'b0;
    437: acceptStates = 1'b0;
    438: acceptStates = 1'b0;
    439: acceptStates = 1'b0;
    440: acceptStates = 1'b0;
    441: acceptStates = 1'b0;
    442: acceptStates = 1'b0;
    443: acceptStates = 1'b0;
    444: acceptStates = 1'b0;
    445: acceptStates = 1'b0;
    446: acceptStates = 1'b0;
    447: acceptStates = 1'b0;
    448: acceptStates = 1'b0;
    449: acceptStates = 1'b0;
    450: acceptStates = 1'b0;
    451: acceptStates = 1'b0;
    452: acceptStates = 1'b0;
    453: acceptStates = 1'b0;
    454: acceptStates = 1'b0;
    455: acceptStates = 1'b0;
    456: acceptStates = 1'b0;
    457: acceptStates = 1'b0;
    458: acceptStates = 1'b0;
    459: acceptStates = 1'b0;
    460: acceptStates = 1'b0;
    461: acceptStates = 1'b0;
    462: acceptStates = 1'b0;
    463: acceptStates = 1'b0;
    464: acceptStates = 1'b0;
    465: acceptStates = 1'b0;
    466: acceptStates = 1'b0;
    467: acceptStates = 1'b0;
    468: acceptStates = 1'b0;
    469: acceptStates = 1'b0;
    470: acceptStates = 1'b0;
    471: acceptStates = 1'b0;
    472: acceptStates = 1'b0;
    473: acceptStates = 1'b0;
    474: acceptStates = 1'b0;
    475: acceptStates = 1'b0;
    476: acceptStates = 1'b0;
    477: acceptStates = 1'b0;
    478: acceptStates = 1'b0;
    479: acceptStates = 1'b0;
    480: acceptStates = 1'b0;
    481: acceptStates = 1'b0;
    482: acceptStates = 1'b0;
    483: acceptStates = 1'b0;
    484: acceptStates = 1'b0;
    485: acceptStates = 1'b0;
    486: acceptStates = 1'b0;
    487: acceptStates = 1'b0;
    488: acceptStates = 1'b0;
    489: acceptStates = 1'b0;
    490: acceptStates = 1'b0;
    491: acceptStates = 1'b0;
    492: acceptStates = 1'b0;
    493: acceptStates = 1'b0;
    494: acceptStates = 1'b0;
    495: acceptStates = 1'b0;
    496: acceptStates = 1'b0;
    497: acceptStates = 1'b0;
    498: acceptStates = 1'b0;
    499: acceptStates = 1'b0;
    500: acceptStates = 1'b0;
    501: acceptStates = 1'b0;
    502: acceptStates = 1'b0;
    503: acceptStates = 1'b0;
    504: acceptStates = 1'b0;
    505: acceptStates = 1'b0;
    506: acceptStates = 1'b0;
    507: acceptStates = 1'b0;
    508: acceptStates = 1'b0;
    509: acceptStates = 1'b0;
    510: acceptStates = 1'b0;
    511: acceptStates = 1'b0;
    512: acceptStates = 1'b0;
    513: acceptStates = 1'b0;
    514: acceptStates = 1'b0;
    515: acceptStates = 1'b0;
    516: acceptStates = 1'b0;
    517: acceptStates = 1'b0;
    518: acceptStates = 1'b0;
    519: acceptStates = 1'b0;
    520: acceptStates = 1'b0;
    521: acceptStates = 1'b0;
    522: acceptStates = 1'b0;
    523: acceptStates = 1'b0;
    524: acceptStates = 1'b0;
    525: acceptStates = 1'b0;
    526: acceptStates = 1'b0;
    527: acceptStates = 1'b0;
    528: acceptStates = 1'b0;
    529: acceptStates = 1'b0;
    530: acceptStates = 1'b0;
    531: acceptStates = 1'b0;
    532: acceptStates = 1'b0;
    533: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd1;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd6;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd7;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd8;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd9;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd10;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd12;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd13;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd14;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd15;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd16;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd16;
      12: stateTransition = 11'd16;
      13: stateTransition = 11'd17;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd18;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd20;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd21;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd22;
      12: stateTransition = 11'd22;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd533;
      2: stateTransition = 11'd533;
      3: stateTransition = 11'd533;
      4: stateTransition = 11'd533;
      5: stateTransition = 11'd533;
      6: stateTransition = 11'd533;
      7: stateTransition = 11'd533;
      8: stateTransition = 11'd533;
      9: stateTransition = 11'd533;
      10: stateTransition = 11'd533;
      11: stateTransition = 11'd533;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd533;
      14: stateTransition = 11'd533;
      15: stateTransition = 11'd533;
      16: stateTransition = 11'd533;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd2;
      2: stateTransition = 11'd2;
      3: stateTransition = 11'd2;
      4: stateTransition = 11'd2;
      5: stateTransition = 11'd2;
      6: stateTransition = 11'd2;
      7: stateTransition = 11'd2;
      8: stateTransition = 11'd2;
      9: stateTransition = 11'd2;
      10: stateTransition = 11'd2;
      11: stateTransition = 11'd2;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd2;
      14: stateTransition = 11'd2;
      15: stateTransition = 11'd2;
      16: stateTransition = 11'd2;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd23;
      2: stateTransition = 11'd23;
      3: stateTransition = 11'd23;
      4: stateTransition = 11'd23;
      5: stateTransition = 11'd23;
      6: stateTransition = 11'd23;
      7: stateTransition = 11'd23;
      8: stateTransition = 11'd23;
      9: stateTransition = 11'd23;
      10: stateTransition = 11'd23;
      11: stateTransition = 11'd23;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd23;
      14: stateTransition = 11'd23;
      15: stateTransition = 11'd23;
      16: stateTransition = 11'd23;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd24;
      5: stateTransition = 11'd24;
      6: stateTransition = 11'd24;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd24;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd25;
      2: stateTransition = 11'd25;
      3: stateTransition = 11'd25;
      4: stateTransition = 11'd25;
      5: stateTransition = 11'd25;
      6: stateTransition = 11'd25;
      7: stateTransition = 11'd25;
      8: stateTransition = 11'd25;
      9: stateTransition = 11'd25;
      10: stateTransition = 11'd25;
      11: stateTransition = 11'd25;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd25;
      14: stateTransition = 11'd25;
      15: stateTransition = 11'd25;
      16: stateTransition = 11'd25;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd26;
      2: stateTransition = 11'd26;
      3: stateTransition = 11'd26;
      4: stateTransition = 11'd26;
      5: stateTransition = 11'd26;
      6: stateTransition = 11'd26;
      7: stateTransition = 11'd26;
      8: stateTransition = 11'd26;
      9: stateTransition = 11'd26;
      10: stateTransition = 11'd26;
      11: stateTransition = 11'd26;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd26;
      14: stateTransition = 11'd26;
      15: stateTransition = 11'd26;
      16: stateTransition = 11'd26;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd28;
      2: stateTransition = 11'd28;
      3: stateTransition = 11'd28;
      4: stateTransition = 11'd28;
      5: stateTransition = 11'd28;
      6: stateTransition = 11'd28;
      7: stateTransition = 11'd28;
      8: stateTransition = 11'd28;
      9: stateTransition = 11'd28;
      10: stateTransition = 11'd28;
      11: stateTransition = 11'd28;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd28;
      14: stateTransition = 11'd28;
      15: stateTransition = 11'd28;
      16: stateTransition = 11'd28;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd29;
      2: stateTransition = 11'd29;
      3: stateTransition = 11'd29;
      4: stateTransition = 11'd29;
      5: stateTransition = 11'd29;
      6: stateTransition = 11'd29;
      7: stateTransition = 11'd29;
      8: stateTransition = 11'd29;
      9: stateTransition = 11'd29;
      10: stateTransition = 11'd29;
      11: stateTransition = 11'd29;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd29;
      14: stateTransition = 11'd29;
      15: stateTransition = 11'd29;
      16: stateTransition = 11'd29;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd30;
      3: stateTransition = 11'd30;
      4: stateTransition = 11'd30;
      5: stateTransition = 11'd30;
      6: stateTransition = 11'd30;
      7: stateTransition = 11'd30;
      8: stateTransition = 11'd30;
      9: stateTransition = 11'd30;
      10: stateTransition = 11'd30;
      11: stateTransition = 11'd30;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd30;
      14: stateTransition = 11'd30;
      15: stateTransition = 11'd30;
      16: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd31;
      2: stateTransition = 11'd31;
      3: stateTransition = 11'd31;
      4: stateTransition = 11'd31;
      5: stateTransition = 11'd31;
      6: stateTransition = 11'd31;
      7: stateTransition = 11'd31;
      8: stateTransition = 11'd31;
      9: stateTransition = 11'd31;
      10: stateTransition = 11'd31;
      11: stateTransition = 11'd31;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd31;
      14: stateTransition = 11'd31;
      15: stateTransition = 11'd31;
      16: stateTransition = 11'd31;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd32;
      2: stateTransition = 11'd32;
      3: stateTransition = 11'd32;
      4: stateTransition = 11'd32;
      5: stateTransition = 11'd32;
      6: stateTransition = 11'd32;
      7: stateTransition = 11'd32;
      8: stateTransition = 11'd32;
      9: stateTransition = 11'd32;
      10: stateTransition = 11'd32;
      11: stateTransition = 11'd32;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd32;
      14: stateTransition = 11'd32;
      15: stateTransition = 11'd32;
      16: stateTransition = 11'd32;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd33;
      2: stateTransition = 11'd33;
      3: stateTransition = 11'd33;
      4: stateTransition = 11'd33;
      5: stateTransition = 11'd33;
      6: stateTransition = 11'd33;
      7: stateTransition = 11'd33;
      8: stateTransition = 11'd33;
      9: stateTransition = 11'd33;
      10: stateTransition = 11'd33;
      11: stateTransition = 11'd33;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd33;
      14: stateTransition = 11'd33;
      15: stateTransition = 11'd33;
      16: stateTransition = 11'd33;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd34;
      2: stateTransition = 11'd34;
      3: stateTransition = 11'd34;
      4: stateTransition = 11'd34;
      5: stateTransition = 11'd34;
      6: stateTransition = 11'd34;
      7: stateTransition = 11'd34;
      8: stateTransition = 11'd34;
      9: stateTransition = 11'd34;
      10: stateTransition = 11'd34;
      11: stateTransition = 11'd34;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd34;
      14: stateTransition = 11'd34;
      15: stateTransition = 11'd34;
      16: stateTransition = 11'd34;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd35;
      2: stateTransition = 11'd35;
      3: stateTransition = 11'd35;
      4: stateTransition = 11'd35;
      5: stateTransition = 11'd35;
      6: stateTransition = 11'd35;
      7: stateTransition = 11'd35;
      8: stateTransition = 11'd35;
      9: stateTransition = 11'd35;
      10: stateTransition = 11'd35;
      11: stateTransition = 11'd35;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd35;
      14: stateTransition = 11'd35;
      15: stateTransition = 11'd35;
      16: stateTransition = 11'd35;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd36;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd36;
      4: stateTransition = 11'd36;
      5: stateTransition = 11'd36;
      6: stateTransition = 11'd36;
      7: stateTransition = 11'd36;
      8: stateTransition = 11'd36;
      9: stateTransition = 11'd36;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd36;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd36;
      14: stateTransition = 11'd36;
      15: stateTransition = 11'd36;
      16: stateTransition = 11'd36;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd37;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd37;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd37;
      6: stateTransition = 11'd37;
      7: stateTransition = 11'd37;
      8: stateTransition = 11'd37;
      9: stateTransition = 11'd37;
      10: stateTransition = 11'd37;
      11: stateTransition = 11'd37;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd37;
      14: stateTransition = 11'd37;
      15: stateTransition = 11'd37;
      16: stateTransition = 11'd37;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd38;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd38;
      4: stateTransition = 11'd38;
      5: stateTransition = 11'd38;
      6: stateTransition = 11'd38;
      7: stateTransition = 11'd38;
      8: stateTransition = 11'd38;
      9: stateTransition = 11'd38;
      10: stateTransition = 11'd38;
      11: stateTransition = 11'd38;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd38;
      14: stateTransition = 11'd38;
      15: stateTransition = 11'd38;
      16: stateTransition = 11'd38;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd39;
      2: stateTransition = 11'd39;
      3: stateTransition = 11'd39;
      4: stateTransition = 11'd39;
      5: stateTransition = 11'd39;
      6: stateTransition = 11'd39;
      7: stateTransition = 11'd39;
      8: stateTransition = 11'd39;
      9: stateTransition = 11'd39;
      10: stateTransition = 11'd39;
      11: stateTransition = 11'd39;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd39;
      14: stateTransition = 11'd39;
      15: stateTransition = 11'd39;
      16: stateTransition = 11'd39;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd40;
      2: stateTransition = 11'd40;
      3: stateTransition = 11'd40;
      4: stateTransition = 11'd40;
      5: stateTransition = 11'd40;
      6: stateTransition = 11'd40;
      7: stateTransition = 11'd40;
      8: stateTransition = 11'd40;
      9: stateTransition = 11'd40;
      10: stateTransition = 11'd40;
      11: stateTransition = 11'd40;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd40;
      14: stateTransition = 11'd40;
      15: stateTransition = 11'd40;
      16: stateTransition = 11'd40;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd41;
      2: stateTransition = 11'd41;
      3: stateTransition = 11'd41;
      4: stateTransition = 11'd41;
      5: stateTransition = 11'd41;
      6: stateTransition = 11'd41;
      7: stateTransition = 11'd41;
      8: stateTransition = 11'd41;
      9: stateTransition = 11'd41;
      10: stateTransition = 11'd41;
      11: stateTransition = 11'd41;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd41;
      14: stateTransition = 11'd41;
      15: stateTransition = 11'd41;
      16: stateTransition = 11'd41;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd42;
      2: stateTransition = 11'd42;
      3: stateTransition = 11'd42;
      4: stateTransition = 11'd42;
      5: stateTransition = 11'd42;
      6: stateTransition = 11'd42;
      7: stateTransition = 11'd42;
      8: stateTransition = 11'd42;
      9: stateTransition = 11'd42;
      10: stateTransition = 11'd42;
      11: stateTransition = 11'd42;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd42;
      14: stateTransition = 11'd42;
      15: stateTransition = 11'd42;
      16: stateTransition = 11'd42;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd43;
      2: stateTransition = 11'd43;
      3: stateTransition = 11'd43;
      4: stateTransition = 11'd43;
      5: stateTransition = 11'd43;
      6: stateTransition = 11'd43;
      7: stateTransition = 11'd43;
      8: stateTransition = 11'd43;
      9: stateTransition = 11'd43;
      10: stateTransition = 11'd43;
      11: stateTransition = 11'd43;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd43;
      14: stateTransition = 11'd43;
      15: stateTransition = 11'd43;
      16: stateTransition = 11'd43;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd44;
      2: stateTransition = 11'd44;
      3: stateTransition = 11'd44;
      4: stateTransition = 11'd44;
      5: stateTransition = 11'd44;
      6: stateTransition = 11'd44;
      7: stateTransition = 11'd44;
      8: stateTransition = 11'd44;
      9: stateTransition = 11'd44;
      10: stateTransition = 11'd44;
      11: stateTransition = 11'd44;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd44;
      14: stateTransition = 11'd44;
      15: stateTransition = 11'd44;
      16: stateTransition = 11'd44;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd45;
      2: stateTransition = 11'd45;
      3: stateTransition = 11'd45;
      4: stateTransition = 11'd45;
      5: stateTransition = 11'd45;
      6: stateTransition = 11'd45;
      7: stateTransition = 11'd45;
      8: stateTransition = 11'd45;
      9: stateTransition = 11'd45;
      10: stateTransition = 11'd45;
      11: stateTransition = 11'd45;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd45;
      14: stateTransition = 11'd45;
      15: stateTransition = 11'd45;
      16: stateTransition = 11'd45;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd46;
      2: stateTransition = 11'd46;
      3: stateTransition = 11'd46;
      4: stateTransition = 11'd46;
      5: stateTransition = 11'd46;
      6: stateTransition = 11'd46;
      7: stateTransition = 11'd46;
      8: stateTransition = 11'd46;
      9: stateTransition = 11'd46;
      10: stateTransition = 11'd46;
      11: stateTransition = 11'd46;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd46;
      14: stateTransition = 11'd46;
      15: stateTransition = 11'd46;
      16: stateTransition = 11'd46;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd47;
      2: stateTransition = 11'd47;
      3: stateTransition = 11'd47;
      4: stateTransition = 11'd47;
      5: stateTransition = 11'd47;
      6: stateTransition = 11'd47;
      7: stateTransition = 11'd47;
      8: stateTransition = 11'd47;
      9: stateTransition = 11'd47;
      10: stateTransition = 11'd47;
      11: stateTransition = 11'd47;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd47;
      14: stateTransition = 11'd47;
      15: stateTransition = 11'd47;
      16: stateTransition = 11'd47;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd48;
      2: stateTransition = 11'd48;
      3: stateTransition = 11'd48;
      4: stateTransition = 11'd48;
      5: stateTransition = 11'd48;
      6: stateTransition = 11'd48;
      7: stateTransition = 11'd48;
      8: stateTransition = 11'd48;
      9: stateTransition = 11'd48;
      10: stateTransition = 11'd48;
      11: stateTransition = 11'd48;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd48;
      14: stateTransition = 11'd48;
      15: stateTransition = 11'd48;
      16: stateTransition = 11'd48;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd49;
      2: stateTransition = 11'd49;
      3: stateTransition = 11'd49;
      4: stateTransition = 11'd49;
      5: stateTransition = 11'd49;
      6: stateTransition = 11'd49;
      7: stateTransition = 11'd49;
      8: stateTransition = 11'd49;
      9: stateTransition = 11'd49;
      10: stateTransition = 11'd49;
      11: stateTransition = 11'd49;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd49;
      14: stateTransition = 11'd49;
      15: stateTransition = 11'd49;
      16: stateTransition = 11'd49;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd50;
      2: stateTransition = 11'd50;
      3: stateTransition = 11'd50;
      4: stateTransition = 11'd50;
      5: stateTransition = 11'd50;
      6: stateTransition = 11'd50;
      7: stateTransition = 11'd50;
      8: stateTransition = 11'd50;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd50;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd50;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd51;
      2: stateTransition = 11'd51;
      3: stateTransition = 11'd51;
      4: stateTransition = 11'd51;
      5: stateTransition = 11'd51;
      6: stateTransition = 11'd51;
      7: stateTransition = 11'd51;
      8: stateTransition = 11'd51;
      9: stateTransition = 11'd51;
      10: stateTransition = 11'd51;
      11: stateTransition = 11'd51;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd51;
      14: stateTransition = 11'd51;
      15: stateTransition = 11'd51;
      16: stateTransition = 11'd51;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd52;
      3: stateTransition = 11'd52;
      4: stateTransition = 11'd52;
      5: stateTransition = 11'd52;
      6: stateTransition = 11'd52;
      7: stateTransition = 11'd52;
      8: stateTransition = 11'd52;
      9: stateTransition = 11'd52;
      10: stateTransition = 11'd52;
      11: stateTransition = 11'd52;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd52;
      14: stateTransition = 11'd52;
      15: stateTransition = 11'd52;
      16: stateTransition = 11'd52;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd53;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd53;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd53;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd54;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd54;
      4: stateTransition = 11'd54;
      5: stateTransition = 11'd54;
      6: stateTransition = 11'd54;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd54;
      10: stateTransition = 11'd54;
      11: stateTransition = 11'd54;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd54;
      14: stateTransition = 11'd54;
      15: stateTransition = 11'd54;
      16: stateTransition = 11'd54;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd55;
      2: stateTransition = 11'd55;
      3: stateTransition = 11'd55;
      4: stateTransition = 11'd55;
      5: stateTransition = 11'd55;
      6: stateTransition = 11'd55;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd55;
      10: stateTransition = 11'd55;
      11: stateTransition = 11'd55;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd55;
      14: stateTransition = 11'd55;
      15: stateTransition = 11'd55;
      16: stateTransition = 11'd55;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd56;
      2: stateTransition = 11'd56;
      3: stateTransition = 11'd56;
      4: stateTransition = 11'd56;
      5: stateTransition = 11'd56;
      6: stateTransition = 11'd56;
      7: stateTransition = 11'd56;
      8: stateTransition = 11'd56;
      9: stateTransition = 11'd56;
      10: stateTransition = 11'd56;
      11: stateTransition = 11'd56;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd56;
      14: stateTransition = 11'd56;
      15: stateTransition = 11'd56;
      16: stateTransition = 11'd56;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd57;
      2: stateTransition = 11'd57;
      3: stateTransition = 11'd57;
      4: stateTransition = 11'd57;
      5: stateTransition = 11'd57;
      6: stateTransition = 11'd57;
      7: stateTransition = 11'd57;
      8: stateTransition = 11'd57;
      9: stateTransition = 11'd57;
      10: stateTransition = 11'd57;
      11: stateTransition = 11'd57;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd57;
      14: stateTransition = 11'd57;
      15: stateTransition = 11'd57;
      16: stateTransition = 11'd57;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd58;
      3: stateTransition = 11'd58;
      4: stateTransition = 11'd58;
      5: stateTransition = 11'd58;
      6: stateTransition = 11'd58;
      7: stateTransition = 11'd58;
      8: stateTransition = 11'd58;
      9: stateTransition = 11'd58;
      10: stateTransition = 11'd58;
      11: stateTransition = 11'd58;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd58;
      14: stateTransition = 11'd58;
      15: stateTransition = 11'd58;
      16: stateTransition = 11'd58;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd59;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd59;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd59;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    60: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd60;
      2: stateTransition = 11'd60;
      3: stateTransition = 11'd60;
      4: stateTransition = 11'd60;
      5: stateTransition = 11'd60;
      6: stateTransition = 11'd60;
      7: stateTransition = 11'd60;
      8: stateTransition = 11'd60;
      9: stateTransition = 11'd60;
      10: stateTransition = 11'd60;
      11: stateTransition = 11'd60;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd60;
      14: stateTransition = 11'd60;
      15: stateTransition = 11'd60;
      16: stateTransition = 11'd60;
      default: stateTransition = 11'bX;
    endcase
    61: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd61;
      2: stateTransition = 11'd61;
      3: stateTransition = 11'd61;
      4: stateTransition = 11'd61;
      5: stateTransition = 11'd61;
      6: stateTransition = 11'd61;
      7: stateTransition = 11'd61;
      8: stateTransition = 11'd61;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd61;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd61;
      default: stateTransition = 11'bX;
    endcase
    62: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd62;
      2: stateTransition = 11'd62;
      3: stateTransition = 11'd62;
      4: stateTransition = 11'd62;
      5: stateTransition = 11'd62;
      6: stateTransition = 11'd62;
      7: stateTransition = 11'd62;
      8: stateTransition = 11'd62;
      9: stateTransition = 11'd62;
      10: stateTransition = 11'd62;
      11: stateTransition = 11'd62;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd62;
      14: stateTransition = 11'd62;
      15: stateTransition = 11'd62;
      16: stateTransition = 11'd62;
      default: stateTransition = 11'bX;
    endcase
    63: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd63;
      2: stateTransition = 11'd63;
      3: stateTransition = 11'd63;
      4: stateTransition = 11'd63;
      5: stateTransition = 11'd63;
      6: stateTransition = 11'd63;
      7: stateTransition = 11'd63;
      8: stateTransition = 11'd63;
      9: stateTransition = 11'd63;
      10: stateTransition = 11'd63;
      11: stateTransition = 11'd63;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd63;
      14: stateTransition = 11'd63;
      15: stateTransition = 11'd63;
      16: stateTransition = 11'd63;
      default: stateTransition = 11'bX;
    endcase
    64: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd64;
      5: stateTransition = 11'd64;
      6: stateTransition = 11'd64;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    65: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd65;
      2: stateTransition = 11'd65;
      3: stateTransition = 11'd65;
      4: stateTransition = 11'd65;
      5: stateTransition = 11'd65;
      6: stateTransition = 11'd65;
      7: stateTransition = 11'd65;
      8: stateTransition = 11'd65;
      9: stateTransition = 11'd65;
      10: stateTransition = 11'd65;
      11: stateTransition = 11'd65;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd65;
      14: stateTransition = 11'd65;
      15: stateTransition = 11'd65;
      16: stateTransition = 11'd65;
      default: stateTransition = 11'bX;
    endcase
    66: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd66;
      2: stateTransition = 11'd66;
      3: stateTransition = 11'd66;
      4: stateTransition = 11'd66;
      5: stateTransition = 11'd66;
      6: stateTransition = 11'd66;
      7: stateTransition = 11'd66;
      8: stateTransition = 11'd66;
      9: stateTransition = 11'd66;
      10: stateTransition = 11'd66;
      11: stateTransition = 11'd66;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd66;
      14: stateTransition = 11'd66;
      15: stateTransition = 11'd66;
      16: stateTransition = 11'd66;
      default: stateTransition = 11'bX;
    endcase
    67: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd67;
      2: stateTransition = 11'd67;
      3: stateTransition = 11'd67;
      4: stateTransition = 11'd67;
      5: stateTransition = 11'd67;
      6: stateTransition = 11'd67;
      7: stateTransition = 11'd67;
      8: stateTransition = 11'd67;
      9: stateTransition = 11'd67;
      10: stateTransition = 11'd67;
      11: stateTransition = 11'd67;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd67;
      14: stateTransition = 11'd67;
      15: stateTransition = 11'd67;
      16: stateTransition = 11'd67;
      default: stateTransition = 11'bX;
    endcase
    68: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd68;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd68;
      4: stateTransition = 11'd68;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd68;
      7: stateTransition = 11'd68;
      8: stateTransition = 11'd68;
      9: stateTransition = 11'd68;
      10: stateTransition = 11'd68;
      11: stateTransition = 11'd68;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd68;
      14: stateTransition = 11'd68;
      15: stateTransition = 11'd68;
      16: stateTransition = 11'd68;
      default: stateTransition = 11'bX;
    endcase
    69: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd69;
      2: stateTransition = 11'd69;
      3: stateTransition = 11'd69;
      4: stateTransition = 11'd69;
      5: stateTransition = 11'd69;
      6: stateTransition = 11'd69;
      7: stateTransition = 11'd69;
      8: stateTransition = 11'd69;
      9: stateTransition = 11'd69;
      10: stateTransition = 11'd69;
      11: stateTransition = 11'd69;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd69;
      14: stateTransition = 11'd69;
      15: stateTransition = 11'd69;
      16: stateTransition = 11'd69;
      default: stateTransition = 11'bX;
    endcase
    70: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd70;
      2: stateTransition = 11'd70;
      3: stateTransition = 11'd70;
      4: stateTransition = 11'd70;
      5: stateTransition = 11'd70;
      6: stateTransition = 11'd70;
      7: stateTransition = 11'd70;
      8: stateTransition = 11'd70;
      9: stateTransition = 11'd70;
      10: stateTransition = 11'd70;
      11: stateTransition = 11'd70;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd70;
      14: stateTransition = 11'd70;
      15: stateTransition = 11'd70;
      16: stateTransition = 11'd70;
      default: stateTransition = 11'bX;
    endcase
    71: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd71;
      2: stateTransition = 11'd71;
      3: stateTransition = 11'd71;
      4: stateTransition = 11'd71;
      5: stateTransition = 11'd71;
      6: stateTransition = 11'd71;
      7: stateTransition = 11'd71;
      8: stateTransition = 11'd71;
      9: stateTransition = 11'd71;
      10: stateTransition = 11'd71;
      11: stateTransition = 11'd71;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd71;
      14: stateTransition = 11'd71;
      15: stateTransition = 11'd71;
      16: stateTransition = 11'd71;
      default: stateTransition = 11'bX;
    endcase
    72: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd72;
      2: stateTransition = 11'd72;
      3: stateTransition = 11'd72;
      4: stateTransition = 11'd72;
      5: stateTransition = 11'd72;
      6: stateTransition = 11'd72;
      7: stateTransition = 11'd72;
      8: stateTransition = 11'd72;
      9: stateTransition = 11'd72;
      10: stateTransition = 11'd72;
      11: stateTransition = 11'd72;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd72;
      14: stateTransition = 11'd72;
      15: stateTransition = 11'd72;
      16: stateTransition = 11'd72;
      default: stateTransition = 11'bX;
    endcase
    73: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd73;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd73;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd73;
      8: stateTransition = 11'd73;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      default: stateTransition = 11'bX;
    endcase
    74: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd74;
      2: stateTransition = 11'd74;
      3: stateTransition = 11'd74;
      4: stateTransition = 11'd74;
      5: stateTransition = 11'd74;
      6: stateTransition = 11'd74;
      7: stateTransition = 11'd74;
      8: stateTransition = 11'd74;
      9: stateTransition = 11'd74;
      10: stateTransition = 11'd74;
      11: stateTransition = 11'd74;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd74;
      14: stateTransition = 11'd74;
      15: stateTransition = 11'd74;
      16: stateTransition = 11'd74;
      default: stateTransition = 11'bX;
    endcase
    75: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd75;
      2: stateTransition = 11'd75;
      3: stateTransition = 11'd75;
      4: stateTransition = 11'd75;
      5: stateTransition = 11'd75;
      6: stateTransition = 11'd75;
      7: stateTransition = 11'd75;
      8: stateTransition = 11'd75;
      9: stateTransition = 11'd75;
      10: stateTransition = 11'd75;
      11: stateTransition = 11'd75;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd75;
      14: stateTransition = 11'd75;
      15: stateTransition = 11'd75;
      16: stateTransition = 11'd75;
      default: stateTransition = 11'bX;
    endcase
    76: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd76;
      2: stateTransition = 11'd76;
      3: stateTransition = 11'd76;
      4: stateTransition = 11'd76;
      5: stateTransition = 11'd76;
      6: stateTransition = 11'd76;
      7: stateTransition = 11'd76;
      8: stateTransition = 11'd76;
      9: stateTransition = 11'd76;
      10: stateTransition = 11'd76;
      11: stateTransition = 11'd76;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd76;
      14: stateTransition = 11'd76;
      15: stateTransition = 11'd76;
      16: stateTransition = 11'd76;
      default: stateTransition = 11'bX;
    endcase
    77: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd77;
      2: stateTransition = 11'd77;
      3: stateTransition = 11'd77;
      4: stateTransition = 11'd77;
      5: stateTransition = 11'd77;
      6: stateTransition = 11'd77;
      7: stateTransition = 11'd77;
      8: stateTransition = 11'd77;
      9: stateTransition = 11'd77;
      10: stateTransition = 11'd77;
      11: stateTransition = 11'd77;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd77;
      14: stateTransition = 11'd77;
      15: stateTransition = 11'd77;
      16: stateTransition = 11'd77;
      default: stateTransition = 11'bX;
    endcase
    78: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd78;
      2: stateTransition = 11'd78;
      3: stateTransition = 11'd78;
      4: stateTransition = 11'd78;
      5: stateTransition = 11'd78;
      6: stateTransition = 11'd78;
      7: stateTransition = 11'd78;
      8: stateTransition = 11'd78;
      9: stateTransition = 11'd78;
      10: stateTransition = 11'd78;
      11: stateTransition = 11'd78;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd78;
      14: stateTransition = 11'd78;
      15: stateTransition = 11'd78;
      16: stateTransition = 11'd78;
      default: stateTransition = 11'bX;
    endcase
    79: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd79;
      2: stateTransition = 11'd79;
      3: stateTransition = 11'd79;
      4: stateTransition = 11'd79;
      5: stateTransition = 11'd79;
      6: stateTransition = 11'd79;
      7: stateTransition = 11'd79;
      8: stateTransition = 11'd79;
      9: stateTransition = 11'd79;
      10: stateTransition = 11'd79;
      11: stateTransition = 11'd79;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd79;
      14: stateTransition = 11'd79;
      15: stateTransition = 11'd79;
      16: stateTransition = 11'd79;
      default: stateTransition = 11'bX;
    endcase
    80: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd80;
      2: stateTransition = 11'd80;
      3: stateTransition = 11'd80;
      4: stateTransition = 11'd80;
      5: stateTransition = 11'd80;
      6: stateTransition = 11'd80;
      7: stateTransition = 11'd80;
      8: stateTransition = 11'd80;
      9: stateTransition = 11'd80;
      10: stateTransition = 11'd80;
      11: stateTransition = 11'd80;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd80;
      14: stateTransition = 11'd80;
      15: stateTransition = 11'd80;
      16: stateTransition = 11'd80;
      default: stateTransition = 11'bX;
    endcase
    81: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd81;
      2: stateTransition = 11'd81;
      3: stateTransition = 11'd81;
      4: stateTransition = 11'd81;
      5: stateTransition = 11'd81;
      6: stateTransition = 11'd81;
      7: stateTransition = 11'd81;
      8: stateTransition = 11'd81;
      9: stateTransition = 11'd81;
      10: stateTransition = 11'd81;
      11: stateTransition = 11'd81;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd81;
      14: stateTransition = 11'd81;
      15: stateTransition = 11'd81;
      16: stateTransition = 11'd81;
      default: stateTransition = 11'bX;
    endcase
    82: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd82;
      2: stateTransition = 11'd82;
      3: stateTransition = 11'd82;
      4: stateTransition = 11'd82;
      5: stateTransition = 11'd82;
      6: stateTransition = 11'd82;
      7: stateTransition = 11'd82;
      8: stateTransition = 11'd82;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd82;
      11: stateTransition = 11'd82;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd82;
      14: stateTransition = 11'd82;
      15: stateTransition = 11'd82;
      16: stateTransition = 11'd82;
      default: stateTransition = 11'bX;
    endcase
    83: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd83;
      2: stateTransition = 11'd83;
      3: stateTransition = 11'd83;
      4: stateTransition = 11'd83;
      5: stateTransition = 11'd83;
      6: stateTransition = 11'd83;
      7: stateTransition = 11'd83;
      8: stateTransition = 11'd83;
      9: stateTransition = 11'd83;
      10: stateTransition = 11'd83;
      11: stateTransition = 11'd83;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd83;
      14: stateTransition = 11'd83;
      15: stateTransition = 11'd83;
      16: stateTransition = 11'd83;
      default: stateTransition = 11'bX;
    endcase
    84: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd84;
      2: stateTransition = 11'd84;
      3: stateTransition = 11'd84;
      4: stateTransition = 11'd84;
      5: stateTransition = 11'd84;
      6: stateTransition = 11'd84;
      7: stateTransition = 11'd84;
      8: stateTransition = 11'd84;
      9: stateTransition = 11'd84;
      10: stateTransition = 11'd84;
      11: stateTransition = 11'd84;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd84;
      14: stateTransition = 11'd84;
      15: stateTransition = 11'd84;
      16: stateTransition = 11'd84;
      default: stateTransition = 11'bX;
    endcase
    85: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd85;
      2: stateTransition = 11'd85;
      3: stateTransition = 11'd85;
      4: stateTransition = 11'd85;
      5: stateTransition = 11'd85;
      6: stateTransition = 11'd85;
      7: stateTransition = 11'd85;
      8: stateTransition = 11'd85;
      9: stateTransition = 11'd85;
      10: stateTransition = 11'd85;
      11: stateTransition = 11'd85;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd85;
      14: stateTransition = 11'd85;
      15: stateTransition = 11'd85;
      16: stateTransition = 11'd85;
      default: stateTransition = 11'bX;
    endcase
    86: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd86;
      2: stateTransition = 11'd86;
      3: stateTransition = 11'd86;
      4: stateTransition = 11'd86;
      5: stateTransition = 11'd86;
      6: stateTransition = 11'd86;
      7: stateTransition = 11'd86;
      8: stateTransition = 11'd86;
      9: stateTransition = 11'd86;
      10: stateTransition = 11'd86;
      11: stateTransition = 11'd86;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd86;
      14: stateTransition = 11'd86;
      15: stateTransition = 11'd86;
      16: stateTransition = 11'd86;
      default: stateTransition = 11'bX;
    endcase
    87: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd87;
      2: stateTransition = 11'd87;
      3: stateTransition = 11'd87;
      4: stateTransition = 11'd87;
      5: stateTransition = 11'd87;
      6: stateTransition = 11'd87;
      7: stateTransition = 11'd87;
      8: stateTransition = 11'd87;
      9: stateTransition = 11'd87;
      10: stateTransition = 11'd87;
      11: stateTransition = 11'd87;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd87;
      14: stateTransition = 11'd87;
      15: stateTransition = 11'd87;
      16: stateTransition = 11'd87;
      default: stateTransition = 11'bX;
    endcase
    88: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd88;
      2: stateTransition = 11'd88;
      3: stateTransition = 11'd88;
      4: stateTransition = 11'd88;
      5: stateTransition = 11'd88;
      6: stateTransition = 11'd88;
      7: stateTransition = 11'd88;
      8: stateTransition = 11'd88;
      9: stateTransition = 11'd88;
      10: stateTransition = 11'd88;
      11: stateTransition = 11'd88;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd88;
      14: stateTransition = 11'd88;
      15: stateTransition = 11'd88;
      16: stateTransition = 11'd88;
      default: stateTransition = 11'bX;
    endcase
    89: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd89;
      2: stateTransition = 11'd89;
      3: stateTransition = 11'd89;
      4: stateTransition = 11'd89;
      5: stateTransition = 11'd89;
      6: stateTransition = 11'd89;
      7: stateTransition = 11'd89;
      8: stateTransition = 11'd89;
      9: stateTransition = 11'd89;
      10: stateTransition = 11'd89;
      11: stateTransition = 11'd89;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd89;
      14: stateTransition = 11'd89;
      15: stateTransition = 11'd89;
      16: stateTransition = 11'd89;
      default: stateTransition = 11'bX;
    endcase
    90: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd90;
      2: stateTransition = 11'd90;
      3: stateTransition = 11'd90;
      4: stateTransition = 11'd90;
      5: stateTransition = 11'd90;
      6: stateTransition = 11'd90;
      7: stateTransition = 11'd90;
      8: stateTransition = 11'd90;
      9: stateTransition = 11'd90;
      10: stateTransition = 11'd90;
      11: stateTransition = 11'd90;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd90;
      14: stateTransition = 11'd90;
      15: stateTransition = 11'd90;
      16: stateTransition = 11'd90;
      default: stateTransition = 11'bX;
    endcase
    91: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd91;
      2: stateTransition = 11'd91;
      3: stateTransition = 11'd91;
      4: stateTransition = 11'd91;
      5: stateTransition = 11'd91;
      6: stateTransition = 11'd91;
      7: stateTransition = 11'd91;
      8: stateTransition = 11'd91;
      9: stateTransition = 11'd91;
      10: stateTransition = 11'd91;
      11: stateTransition = 11'd91;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd91;
      14: stateTransition = 11'd91;
      15: stateTransition = 11'd91;
      16: stateTransition = 11'd91;
      default: stateTransition = 11'bX;
    endcase
    92: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd92;
      2: stateTransition = 11'd92;
      3: stateTransition = 11'd92;
      4: stateTransition = 11'd92;
      5: stateTransition = 11'd92;
      6: stateTransition = 11'd92;
      7: stateTransition = 11'd92;
      8: stateTransition = 11'd92;
      9: stateTransition = 11'd92;
      10: stateTransition = 11'd92;
      11: stateTransition = 11'd92;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd92;
      14: stateTransition = 11'd92;
      15: stateTransition = 11'd92;
      16: stateTransition = 11'd92;
      default: stateTransition = 11'bX;
    endcase
    93: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd93;
      2: stateTransition = 11'd93;
      3: stateTransition = 11'd93;
      4: stateTransition = 11'd93;
      5: stateTransition = 11'd93;
      6: stateTransition = 11'd93;
      7: stateTransition = 11'd93;
      8: stateTransition = 11'd93;
      9: stateTransition = 11'd93;
      10: stateTransition = 11'd93;
      11: stateTransition = 11'd93;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd93;
      14: stateTransition = 11'd93;
      15: stateTransition = 11'd93;
      16: stateTransition = 11'd93;
      default: stateTransition = 11'bX;
    endcase
    94: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd94;
      2: stateTransition = 11'd94;
      3: stateTransition = 11'd94;
      4: stateTransition = 11'd94;
      5: stateTransition = 11'd94;
      6: stateTransition = 11'd94;
      7: stateTransition = 11'd94;
      8: stateTransition = 11'd94;
      9: stateTransition = 11'd94;
      10: stateTransition = 11'd94;
      11: stateTransition = 11'd94;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd94;
      14: stateTransition = 11'd94;
      15: stateTransition = 11'd94;
      16: stateTransition = 11'd94;
      default: stateTransition = 11'bX;
    endcase
    95: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd95;
      2: stateTransition = 11'd95;
      3: stateTransition = 11'd95;
      4: stateTransition = 11'd95;
      5: stateTransition = 11'd95;
      6: stateTransition = 11'd95;
      7: stateTransition = 11'd95;
      8: stateTransition = 11'd95;
      9: stateTransition = 11'd95;
      10: stateTransition = 11'd95;
      11: stateTransition = 11'd95;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd95;
      14: stateTransition = 11'd95;
      15: stateTransition = 11'd95;
      16: stateTransition = 11'd95;
      default: stateTransition = 11'bX;
    endcase
    96: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd96;
      2: stateTransition = 11'd96;
      3: stateTransition = 11'd96;
      4: stateTransition = 11'd96;
      5: stateTransition = 11'd96;
      6: stateTransition = 11'd96;
      7: stateTransition = 11'd96;
      8: stateTransition = 11'd96;
      9: stateTransition = 11'd96;
      10: stateTransition = 11'd96;
      11: stateTransition = 11'd96;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd96;
      14: stateTransition = 11'd96;
      15: stateTransition = 11'd96;
      16: stateTransition = 11'd96;
      default: stateTransition = 11'bX;
    endcase
    97: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd97;
      2: stateTransition = 11'd97;
      3: stateTransition = 11'd97;
      4: stateTransition = 11'd97;
      5: stateTransition = 11'd97;
      6: stateTransition = 11'd97;
      7: stateTransition = 11'd97;
      8: stateTransition = 11'd97;
      9: stateTransition = 11'd97;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd97;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd97;
      14: stateTransition = 11'd97;
      15: stateTransition = 11'd97;
      16: stateTransition = 11'd97;
      default: stateTransition = 11'bX;
    endcase
    98: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd98;
      2: stateTransition = 11'd98;
      3: stateTransition = 11'd98;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd98;
      6: stateTransition = 11'd98;
      7: stateTransition = 11'd98;
      8: stateTransition = 11'd98;
      9: stateTransition = 11'd98;
      10: stateTransition = 11'd98;
      11: stateTransition = 11'd98;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd98;
      14: stateTransition = 11'd98;
      15: stateTransition = 11'd98;
      16: stateTransition = 11'd98;
      default: stateTransition = 11'bX;
    endcase
    99: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd99;
      2: stateTransition = 11'd99;
      3: stateTransition = 11'd99;
      4: stateTransition = 11'd99;
      5: stateTransition = 11'd99;
      6: stateTransition = 11'd99;
      7: stateTransition = 11'd99;
      8: stateTransition = 11'd99;
      9: stateTransition = 11'd99;
      10: stateTransition = 11'd99;
      11: stateTransition = 11'd99;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd99;
      14: stateTransition = 11'd99;
      15: stateTransition = 11'd99;
      16: stateTransition = 11'd99;
      default: stateTransition = 11'bX;
    endcase
    100: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd100;
      2: stateTransition = 11'd100;
      3: stateTransition = 11'd100;
      4: stateTransition = 11'd100;
      5: stateTransition = 11'd100;
      6: stateTransition = 11'd100;
      7: stateTransition = 11'd100;
      8: stateTransition = 11'd100;
      9: stateTransition = 11'd100;
      10: stateTransition = 11'd100;
      11: stateTransition = 11'd100;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd100;
      14: stateTransition = 11'd100;
      15: stateTransition = 11'd100;
      16: stateTransition = 11'd100;
      default: stateTransition = 11'bX;
    endcase
    101: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd101;
      2: stateTransition = 11'd101;
      3: stateTransition = 11'd101;
      4: stateTransition = 11'd101;
      5: stateTransition = 11'd101;
      6: stateTransition = 11'd101;
      7: stateTransition = 11'd101;
      8: stateTransition = 11'd101;
      9: stateTransition = 11'd101;
      10: stateTransition = 11'd101;
      11: stateTransition = 11'd101;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd101;
      14: stateTransition = 11'd101;
      15: stateTransition = 11'd101;
      16: stateTransition = 11'd101;
      default: stateTransition = 11'bX;
    endcase
    102: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd102;
      2: stateTransition = 11'd102;
      3: stateTransition = 11'd102;
      4: stateTransition = 11'd102;
      5: stateTransition = 11'd102;
      6: stateTransition = 11'd102;
      7: stateTransition = 11'd102;
      8: stateTransition = 11'd102;
      9: stateTransition = 11'd102;
      10: stateTransition = 11'd102;
      11: stateTransition = 11'd102;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd102;
      14: stateTransition = 11'd102;
      15: stateTransition = 11'd102;
      16: stateTransition = 11'd102;
      default: stateTransition = 11'bX;
    endcase
    103: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd103;
      2: stateTransition = 11'd103;
      3: stateTransition = 11'd103;
      4: stateTransition = 11'd103;
      5: stateTransition = 11'd103;
      6: stateTransition = 11'd103;
      7: stateTransition = 11'd103;
      8: stateTransition = 11'd103;
      9: stateTransition = 11'd103;
      10: stateTransition = 11'd103;
      11: stateTransition = 11'd103;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd103;
      14: stateTransition = 11'd103;
      15: stateTransition = 11'd103;
      16: stateTransition = 11'd103;
      default: stateTransition = 11'bX;
    endcase
    104: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd104;
      2: stateTransition = 11'd104;
      3: stateTransition = 11'd104;
      4: stateTransition = 11'd104;
      5: stateTransition = 11'd104;
      6: stateTransition = 11'd104;
      7: stateTransition = 11'd104;
      8: stateTransition = 11'd104;
      9: stateTransition = 11'd104;
      10: stateTransition = 11'd104;
      11: stateTransition = 11'd104;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd104;
      14: stateTransition = 11'd104;
      15: stateTransition = 11'd104;
      16: stateTransition = 11'd104;
      default: stateTransition = 11'bX;
    endcase
    105: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    106: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd106;
      2: stateTransition = 11'd106;
      3: stateTransition = 11'd106;
      4: stateTransition = 11'd106;
      5: stateTransition = 11'd106;
      6: stateTransition = 11'd106;
      7: stateTransition = 11'd106;
      8: stateTransition = 11'd106;
      9: stateTransition = 11'd106;
      10: stateTransition = 11'd106;
      11: stateTransition = 11'd106;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd106;
      14: stateTransition = 11'd106;
      15: stateTransition = 11'd106;
      16: stateTransition = 11'd106;
      default: stateTransition = 11'bX;
    endcase
    107: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd107;
      2: stateTransition = 11'd107;
      3: stateTransition = 11'd107;
      4: stateTransition = 11'd107;
      5: stateTransition = 11'd107;
      6: stateTransition = 11'd107;
      7: stateTransition = 11'd107;
      8: stateTransition = 11'd107;
      9: stateTransition = 11'd107;
      10: stateTransition = 11'd107;
      11: stateTransition = 11'd107;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd107;
      14: stateTransition = 11'd107;
      15: stateTransition = 11'd107;
      16: stateTransition = 11'd107;
      default: stateTransition = 11'bX;
    endcase
    108: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd108;
      2: stateTransition = 11'd108;
      3: stateTransition = 11'd108;
      4: stateTransition = 11'd108;
      5: stateTransition = 11'd108;
      6: stateTransition = 11'd108;
      7: stateTransition = 11'd108;
      8: stateTransition = 11'd108;
      9: stateTransition = 11'd108;
      10: stateTransition = 11'd108;
      11: stateTransition = 11'd108;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd108;
      14: stateTransition = 11'd108;
      15: stateTransition = 11'd108;
      16: stateTransition = 11'd108;
      default: stateTransition = 11'bX;
    endcase
    109: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd109;
      2: stateTransition = 11'd109;
      3: stateTransition = 11'd109;
      4: stateTransition = 11'd109;
      5: stateTransition = 11'd109;
      6: stateTransition = 11'd109;
      7: stateTransition = 11'd109;
      8: stateTransition = 11'd109;
      9: stateTransition = 11'd109;
      10: stateTransition = 11'd109;
      11: stateTransition = 11'd109;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd109;
      14: stateTransition = 11'd109;
      15: stateTransition = 11'd109;
      16: stateTransition = 11'd109;
      default: stateTransition = 11'bX;
    endcase
    110: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd110;
      2: stateTransition = 11'd110;
      3: stateTransition = 11'd110;
      4: stateTransition = 11'd110;
      5: stateTransition = 11'd110;
      6: stateTransition = 11'd110;
      7: stateTransition = 11'd110;
      8: stateTransition = 11'd110;
      9: stateTransition = 11'd110;
      10: stateTransition = 11'd110;
      11: stateTransition = 11'd110;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd110;
      14: stateTransition = 11'd110;
      15: stateTransition = 11'd110;
      16: stateTransition = 11'd110;
      default: stateTransition = 11'bX;
    endcase
    111: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd111;
      2: stateTransition = 11'd111;
      3: stateTransition = 11'd111;
      4: stateTransition = 11'd111;
      5: stateTransition = 11'd111;
      6: stateTransition = 11'd111;
      7: stateTransition = 11'd111;
      8: stateTransition = 11'd111;
      9: stateTransition = 11'd111;
      10: stateTransition = 11'd111;
      11: stateTransition = 11'd111;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd111;
      14: stateTransition = 11'd111;
      15: stateTransition = 11'd111;
      16: stateTransition = 11'd111;
      default: stateTransition = 11'bX;
    endcase
    112: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd112;
      2: stateTransition = 11'd112;
      3: stateTransition = 11'd112;
      4: stateTransition = 11'd112;
      5: stateTransition = 11'd112;
      6: stateTransition = 11'd112;
      7: stateTransition = 11'd112;
      8: stateTransition = 11'd112;
      9: stateTransition = 11'd112;
      10: stateTransition = 11'd112;
      11: stateTransition = 11'd112;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd112;
      14: stateTransition = 11'd112;
      15: stateTransition = 11'd112;
      16: stateTransition = 11'd112;
      default: stateTransition = 11'bX;
    endcase
    113: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd113;
      2: stateTransition = 11'd113;
      3: stateTransition = 11'd113;
      4: stateTransition = 11'd113;
      5: stateTransition = 11'd113;
      6: stateTransition = 11'd113;
      7: stateTransition = 11'd113;
      8: stateTransition = 11'd113;
      9: stateTransition = 11'd113;
      10: stateTransition = 11'd113;
      11: stateTransition = 11'd113;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd113;
      14: stateTransition = 11'd113;
      15: stateTransition = 11'd113;
      16: stateTransition = 11'd113;
      default: stateTransition = 11'bX;
    endcase
    114: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd114;
      2: stateTransition = 11'd114;
      3: stateTransition = 11'd114;
      4: stateTransition = 11'd114;
      5: stateTransition = 11'd114;
      6: stateTransition = 11'd114;
      7: stateTransition = 11'd114;
      8: stateTransition = 11'd114;
      9: stateTransition = 11'd114;
      10: stateTransition = 11'd114;
      11: stateTransition = 11'd114;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd114;
      14: stateTransition = 11'd114;
      15: stateTransition = 11'd114;
      16: stateTransition = 11'd114;
      default: stateTransition = 11'bX;
    endcase
    115: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd115;
      2: stateTransition = 11'd115;
      3: stateTransition = 11'd115;
      4: stateTransition = 11'd115;
      5: stateTransition = 11'd115;
      6: stateTransition = 11'd115;
      7: stateTransition = 11'd115;
      8: stateTransition = 11'd115;
      9: stateTransition = 11'd115;
      10: stateTransition = 11'd115;
      11: stateTransition = 11'd115;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd115;
      14: stateTransition = 11'd115;
      15: stateTransition = 11'd115;
      16: stateTransition = 11'd115;
      default: stateTransition = 11'bX;
    endcase
    116: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd116;
      2: stateTransition = 11'd116;
      3: stateTransition = 11'd116;
      4: stateTransition = 11'd116;
      5: stateTransition = 11'd116;
      6: stateTransition = 11'd116;
      7: stateTransition = 11'd116;
      8: stateTransition = 11'd116;
      9: stateTransition = 11'd116;
      10: stateTransition = 11'd116;
      11: stateTransition = 11'd116;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd116;
      14: stateTransition = 11'd116;
      15: stateTransition = 11'd116;
      16: stateTransition = 11'd116;
      default: stateTransition = 11'bX;
    endcase
    117: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd117;
      2: stateTransition = 11'd117;
      3: stateTransition = 11'd117;
      4: stateTransition = 11'd117;
      5: stateTransition = 11'd117;
      6: stateTransition = 11'd117;
      7: stateTransition = 11'd117;
      8: stateTransition = 11'd117;
      9: stateTransition = 11'd117;
      10: stateTransition = 11'd117;
      11: stateTransition = 11'd117;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd117;
      14: stateTransition = 11'd117;
      15: stateTransition = 11'd117;
      16: stateTransition = 11'd117;
      default: stateTransition = 11'bX;
    endcase
    118: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd118;
      2: stateTransition = 11'd118;
      3: stateTransition = 11'd118;
      4: stateTransition = 11'd118;
      5: stateTransition = 11'd118;
      6: stateTransition = 11'd118;
      7: stateTransition = 11'd118;
      8: stateTransition = 11'd118;
      9: stateTransition = 11'd118;
      10: stateTransition = 11'd118;
      11: stateTransition = 11'd118;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd118;
      14: stateTransition = 11'd118;
      15: stateTransition = 11'd118;
      16: stateTransition = 11'd118;
      default: stateTransition = 11'bX;
    endcase
    119: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd119;
      2: stateTransition = 11'd119;
      3: stateTransition = 11'd119;
      4: stateTransition = 11'd119;
      5: stateTransition = 11'd119;
      6: stateTransition = 11'd119;
      7: stateTransition = 11'd119;
      8: stateTransition = 11'd119;
      9: stateTransition = 11'd119;
      10: stateTransition = 11'd119;
      11: stateTransition = 11'd119;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd119;
      14: stateTransition = 11'd119;
      15: stateTransition = 11'd119;
      16: stateTransition = 11'd119;
      default: stateTransition = 11'bX;
    endcase
    120: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd120;
      2: stateTransition = 11'd120;
      3: stateTransition = 11'd120;
      4: stateTransition = 11'd120;
      5: stateTransition = 11'd120;
      6: stateTransition = 11'd120;
      7: stateTransition = 11'd120;
      8: stateTransition = 11'd120;
      9: stateTransition = 11'd120;
      10: stateTransition = 11'd120;
      11: stateTransition = 11'd120;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd120;
      14: stateTransition = 11'd120;
      15: stateTransition = 11'd120;
      16: stateTransition = 11'd120;
      default: stateTransition = 11'bX;
    endcase
    121: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd121;
      2: stateTransition = 11'd121;
      3: stateTransition = 11'd121;
      4: stateTransition = 11'd121;
      5: stateTransition = 11'd121;
      6: stateTransition = 11'd121;
      7: stateTransition = 11'd121;
      8: stateTransition = 11'd121;
      9: stateTransition = 11'd121;
      10: stateTransition = 11'd121;
      11: stateTransition = 11'd121;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd121;
      14: stateTransition = 11'd121;
      15: stateTransition = 11'd121;
      16: stateTransition = 11'd121;
      default: stateTransition = 11'bX;
    endcase
    122: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd122;
      2: stateTransition = 11'd122;
      3: stateTransition = 11'd122;
      4: stateTransition = 11'd122;
      5: stateTransition = 11'd122;
      6: stateTransition = 11'd122;
      7: stateTransition = 11'd122;
      8: stateTransition = 11'd122;
      9: stateTransition = 11'd122;
      10: stateTransition = 11'd122;
      11: stateTransition = 11'd122;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd122;
      14: stateTransition = 11'd122;
      15: stateTransition = 11'd122;
      16: stateTransition = 11'd122;
      default: stateTransition = 11'bX;
    endcase
    123: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd123;
      2: stateTransition = 11'd123;
      3: stateTransition = 11'd123;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd123;
      6: stateTransition = 11'd123;
      7: stateTransition = 11'd123;
      8: stateTransition = 11'd123;
      9: stateTransition = 11'd123;
      10: stateTransition = 11'd123;
      11: stateTransition = 11'd123;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd123;
      14: stateTransition = 11'd123;
      15: stateTransition = 11'd123;
      16: stateTransition = 11'd123;
      default: stateTransition = 11'bX;
    endcase
    124: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd124;
      2: stateTransition = 11'd124;
      3: stateTransition = 11'd124;
      4: stateTransition = 11'd124;
      5: stateTransition = 11'd124;
      6: stateTransition = 11'd124;
      7: stateTransition = 11'd124;
      8: stateTransition = 11'd124;
      9: stateTransition = 11'd124;
      10: stateTransition = 11'd124;
      11: stateTransition = 11'd124;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd124;
      14: stateTransition = 11'd124;
      15: stateTransition = 11'd124;
      16: stateTransition = 11'd124;
      default: stateTransition = 11'bX;
    endcase
    125: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd125;
      2: stateTransition = 11'd125;
      3: stateTransition = 11'd125;
      4: stateTransition = 11'd125;
      5: stateTransition = 11'd125;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd125;
      8: stateTransition = 11'd125;
      9: stateTransition = 11'd125;
      10: stateTransition = 11'd125;
      11: stateTransition = 11'd125;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd125;
      14: stateTransition = 11'd125;
      15: stateTransition = 11'd125;
      16: stateTransition = 11'd125;
      default: stateTransition = 11'bX;
    endcase
    126: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd126;
      5: stateTransition = 11'd126;
      6: stateTransition = 11'd126;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd126;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    127: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd127;
      2: stateTransition = 11'd127;
      3: stateTransition = 11'd127;
      4: stateTransition = 11'd127;
      5: stateTransition = 11'd127;
      6: stateTransition = 11'd127;
      7: stateTransition = 11'd127;
      8: stateTransition = 11'd127;
      9: stateTransition = 11'd127;
      10: stateTransition = 11'd127;
      11: stateTransition = 11'd127;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd127;
      14: stateTransition = 11'd127;
      15: stateTransition = 11'd127;
      16: stateTransition = 11'd127;
      default: stateTransition = 11'bX;
    endcase
    128: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd128;
      2: stateTransition = 11'd128;
      3: stateTransition = 11'd128;
      4: stateTransition = 11'd128;
      5: stateTransition = 11'd128;
      6: stateTransition = 11'd128;
      7: stateTransition = 11'd128;
      8: stateTransition = 11'd128;
      9: stateTransition = 11'd128;
      10: stateTransition = 11'd128;
      11: stateTransition = 11'd128;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd128;
      14: stateTransition = 11'd128;
      15: stateTransition = 11'd128;
      16: stateTransition = 11'd128;
      default: stateTransition = 11'bX;
    endcase
    129: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd129;
      2: stateTransition = 11'd129;
      3: stateTransition = 11'd129;
      4: stateTransition = 11'd129;
      5: stateTransition = 11'd129;
      6: stateTransition = 11'd129;
      7: stateTransition = 11'd129;
      8: stateTransition = 11'd129;
      9: stateTransition = 11'd129;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd129;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd129;
      14: stateTransition = 11'd129;
      15: stateTransition = 11'd129;
      16: stateTransition = 11'd129;
      default: stateTransition = 11'bX;
    endcase
    130: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd130;
      2: stateTransition = 11'd130;
      3: stateTransition = 11'd130;
      4: stateTransition = 11'd130;
      5: stateTransition = 11'd130;
      6: stateTransition = 11'd130;
      7: stateTransition = 11'd130;
      8: stateTransition = 11'd130;
      9: stateTransition = 11'd130;
      10: stateTransition = 11'd130;
      11: stateTransition = 11'd130;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd130;
      14: stateTransition = 11'd130;
      15: stateTransition = 11'd130;
      16: stateTransition = 11'd130;
      default: stateTransition = 11'bX;
    endcase
    131: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd131;
      2: stateTransition = 11'd131;
      3: stateTransition = 11'd131;
      4: stateTransition = 11'd131;
      5: stateTransition = 11'd131;
      6: stateTransition = 11'd131;
      7: stateTransition = 11'd131;
      8: stateTransition = 11'd131;
      9: stateTransition = 11'd131;
      10: stateTransition = 11'd131;
      11: stateTransition = 11'd131;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd131;
      14: stateTransition = 11'd131;
      15: stateTransition = 11'd131;
      16: stateTransition = 11'd131;
      default: stateTransition = 11'bX;
    endcase
    132: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd132;
      2: stateTransition = 11'd132;
      3: stateTransition = 11'd132;
      4: stateTransition = 11'd132;
      5: stateTransition = 11'd132;
      6: stateTransition = 11'd132;
      7: stateTransition = 11'd132;
      8: stateTransition = 11'd132;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd132;
      11: stateTransition = 11'd132;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd132;
      14: stateTransition = 11'd132;
      15: stateTransition = 11'd132;
      16: stateTransition = 11'd132;
      default: stateTransition = 11'bX;
    endcase
    133: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd133;
      2: stateTransition = 11'd133;
      3: stateTransition = 11'd133;
      4: stateTransition = 11'd133;
      5: stateTransition = 11'd133;
      6: stateTransition = 11'd133;
      7: stateTransition = 11'd133;
      8: stateTransition = 11'd133;
      9: stateTransition = 11'd133;
      10: stateTransition = 11'd133;
      11: stateTransition = 11'd133;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd133;
      14: stateTransition = 11'd133;
      15: stateTransition = 11'd133;
      16: stateTransition = 11'd133;
      default: stateTransition = 11'bX;
    endcase
    134: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd134;
      2: stateTransition = 11'd134;
      3: stateTransition = 11'd134;
      4: stateTransition = 11'd134;
      5: stateTransition = 11'd134;
      6: stateTransition = 11'd134;
      7: stateTransition = 11'd134;
      8: stateTransition = 11'd134;
      9: stateTransition = 11'd134;
      10: stateTransition = 11'd134;
      11: stateTransition = 11'd134;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd134;
      14: stateTransition = 11'd134;
      15: stateTransition = 11'd134;
      16: stateTransition = 11'd134;
      default: stateTransition = 11'bX;
    endcase
    135: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd135;
      2: stateTransition = 11'd135;
      3: stateTransition = 11'd135;
      4: stateTransition = 11'd135;
      5: stateTransition = 11'd135;
      6: stateTransition = 11'd135;
      7: stateTransition = 11'd135;
      8: stateTransition = 11'd135;
      9: stateTransition = 11'd135;
      10: stateTransition = 11'd135;
      11: stateTransition = 11'd135;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd135;
      14: stateTransition = 11'd135;
      15: stateTransition = 11'd135;
      16: stateTransition = 11'd135;
      default: stateTransition = 11'bX;
    endcase
    136: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd136;
      2: stateTransition = 11'd136;
      3: stateTransition = 11'd136;
      4: stateTransition = 11'd136;
      5: stateTransition = 11'd136;
      6: stateTransition = 11'd136;
      7: stateTransition = 11'd136;
      8: stateTransition = 11'd136;
      9: stateTransition = 11'd136;
      10: stateTransition = 11'd136;
      11: stateTransition = 11'd136;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd136;
      14: stateTransition = 11'd136;
      15: stateTransition = 11'd136;
      16: stateTransition = 11'd136;
      default: stateTransition = 11'bX;
    endcase
    137: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd137;
      2: stateTransition = 11'd137;
      3: stateTransition = 11'd137;
      4: stateTransition = 11'd137;
      5: stateTransition = 11'd137;
      6: stateTransition = 11'd137;
      7: stateTransition = 11'd137;
      8: stateTransition = 11'd137;
      9: stateTransition = 11'd137;
      10: stateTransition = 11'd137;
      11: stateTransition = 11'd137;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd137;
      14: stateTransition = 11'd137;
      15: stateTransition = 11'd137;
      16: stateTransition = 11'd137;
      default: stateTransition = 11'bX;
    endcase
    138: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd138;
      2: stateTransition = 11'd138;
      3: stateTransition = 11'd138;
      4: stateTransition = 11'd138;
      5: stateTransition = 11'd138;
      6: stateTransition = 11'd138;
      7: stateTransition = 11'd138;
      8: stateTransition = 11'd138;
      9: stateTransition = 11'd138;
      10: stateTransition = 11'd138;
      11: stateTransition = 11'd138;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd138;
      14: stateTransition = 11'd138;
      15: stateTransition = 11'd138;
      16: stateTransition = 11'd138;
      default: stateTransition = 11'bX;
    endcase
    139: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd139;
      2: stateTransition = 11'd139;
      3: stateTransition = 11'd139;
      4: stateTransition = 11'd139;
      5: stateTransition = 11'd139;
      6: stateTransition = 11'd139;
      7: stateTransition = 11'd139;
      8: stateTransition = 11'd139;
      9: stateTransition = 11'd139;
      10: stateTransition = 11'd139;
      11: stateTransition = 11'd139;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd139;
      14: stateTransition = 11'd139;
      15: stateTransition = 11'd139;
      16: stateTransition = 11'd139;
      default: stateTransition = 11'bX;
    endcase
    140: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd140;
      2: stateTransition = 11'd140;
      3: stateTransition = 11'd140;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd140;
      6: stateTransition = 11'd140;
      7: stateTransition = 11'd140;
      8: stateTransition = 11'd140;
      9: stateTransition = 11'd140;
      10: stateTransition = 11'd140;
      11: stateTransition = 11'd140;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd140;
      14: stateTransition = 11'd140;
      15: stateTransition = 11'd140;
      16: stateTransition = 11'd140;
      default: stateTransition = 11'bX;
    endcase
    141: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd141;
      2: stateTransition = 11'd141;
      3: stateTransition = 11'd141;
      4: stateTransition = 11'd141;
      5: stateTransition = 11'd141;
      6: stateTransition = 11'd141;
      7: stateTransition = 11'd141;
      8: stateTransition = 11'd141;
      9: stateTransition = 11'd141;
      10: stateTransition = 11'd141;
      11: stateTransition = 11'd141;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd141;
      14: stateTransition = 11'd141;
      15: stateTransition = 11'd141;
      16: stateTransition = 11'd141;
      default: stateTransition = 11'bX;
    endcase
    142: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd142;
      2: stateTransition = 11'd142;
      3: stateTransition = 11'd142;
      4: stateTransition = 11'd142;
      5: stateTransition = 11'd142;
      6: stateTransition = 11'd142;
      7: stateTransition = 11'd142;
      8: stateTransition = 11'd142;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd142;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd142;
      default: stateTransition = 11'bX;
    endcase
    143: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd143;
      2: stateTransition = 11'd143;
      3: stateTransition = 11'd143;
      4: stateTransition = 11'd143;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd143;
      7: stateTransition = 11'd143;
      8: stateTransition = 11'd143;
      9: stateTransition = 11'd143;
      10: stateTransition = 11'd143;
      11: stateTransition = 11'd143;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd143;
      14: stateTransition = 11'd143;
      15: stateTransition = 11'd143;
      16: stateTransition = 11'd143;
      default: stateTransition = 11'bX;
    endcase
    144: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd144;
      2: stateTransition = 11'd144;
      3: stateTransition = 11'd144;
      4: stateTransition = 11'd144;
      5: stateTransition = 11'd144;
      6: stateTransition = 11'd144;
      7: stateTransition = 11'd144;
      8: stateTransition = 11'd144;
      9: stateTransition = 11'd144;
      10: stateTransition = 11'd144;
      11: stateTransition = 11'd144;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd144;
      14: stateTransition = 11'd144;
      15: stateTransition = 11'd144;
      16: stateTransition = 11'd144;
      default: stateTransition = 11'bX;
    endcase
    145: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd145;
      2: stateTransition = 11'd145;
      3: stateTransition = 11'd145;
      4: stateTransition = 11'd145;
      5: stateTransition = 11'd145;
      6: stateTransition = 11'd145;
      7: stateTransition = 11'd145;
      8: stateTransition = 11'd145;
      9: stateTransition = 11'd145;
      10: stateTransition = 11'd145;
      11: stateTransition = 11'd145;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd145;
      14: stateTransition = 11'd145;
      15: stateTransition = 11'd145;
      16: stateTransition = 11'd145;
      default: stateTransition = 11'bX;
    endcase
    146: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd146;
      2: stateTransition = 11'd146;
      3: stateTransition = 11'd146;
      4: stateTransition = 11'd146;
      5: stateTransition = 11'd146;
      6: stateTransition = 11'd146;
      7: stateTransition = 11'd146;
      8: stateTransition = 11'd146;
      9: stateTransition = 11'd146;
      10: stateTransition = 11'd146;
      11: stateTransition = 11'd146;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd146;
      14: stateTransition = 11'd146;
      15: stateTransition = 11'd146;
      16: stateTransition = 11'd146;
      default: stateTransition = 11'bX;
    endcase
    147: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd147;
      2: stateTransition = 11'd147;
      3: stateTransition = 11'd147;
      4: stateTransition = 11'd147;
      5: stateTransition = 11'd147;
      6: stateTransition = 11'd147;
      7: stateTransition = 11'd147;
      8: stateTransition = 11'd147;
      9: stateTransition = 11'd147;
      10: stateTransition = 11'd147;
      11: stateTransition = 11'd147;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd147;
      14: stateTransition = 11'd147;
      15: stateTransition = 11'd147;
      16: stateTransition = 11'd147;
      default: stateTransition = 11'bX;
    endcase
    148: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd148;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd148;
      4: stateTransition = 11'd148;
      5: stateTransition = 11'd148;
      6: stateTransition = 11'd148;
      7: stateTransition = 11'd148;
      8: stateTransition = 11'd148;
      9: stateTransition = 11'd148;
      10: stateTransition = 11'd148;
      11: stateTransition = 11'd148;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd148;
      14: stateTransition = 11'd148;
      15: stateTransition = 11'd148;
      16: stateTransition = 11'd148;
      default: stateTransition = 11'bX;
    endcase
    149: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd149;
      2: stateTransition = 11'd149;
      3: stateTransition = 11'd149;
      4: stateTransition = 11'd149;
      5: stateTransition = 11'd149;
      6: stateTransition = 11'd149;
      7: stateTransition = 11'd149;
      8: stateTransition = 11'd149;
      9: stateTransition = 11'd149;
      10: stateTransition = 11'd149;
      11: stateTransition = 11'd149;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd149;
      14: stateTransition = 11'd149;
      15: stateTransition = 11'd149;
      16: stateTransition = 11'd149;
      default: stateTransition = 11'bX;
    endcase
    150: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd150;
      2: stateTransition = 11'd150;
      3: stateTransition = 11'd150;
      4: stateTransition = 11'd150;
      5: stateTransition = 11'd150;
      6: stateTransition = 11'd150;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd150;
      9: stateTransition = 11'd150;
      10: stateTransition = 11'd150;
      11: stateTransition = 11'd150;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd150;
      14: stateTransition = 11'd150;
      15: stateTransition = 11'd150;
      16: stateTransition = 11'd150;
      default: stateTransition = 11'bX;
    endcase
    151: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd151;
      2: stateTransition = 11'd151;
      3: stateTransition = 11'd151;
      4: stateTransition = 11'd151;
      5: stateTransition = 11'd151;
      6: stateTransition = 11'd151;
      7: stateTransition = 11'd151;
      8: stateTransition = 11'd151;
      9: stateTransition = 11'd151;
      10: stateTransition = 11'd151;
      11: stateTransition = 11'd151;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd151;
      14: stateTransition = 11'd151;
      15: stateTransition = 11'd151;
      16: stateTransition = 11'd151;
      default: stateTransition = 11'bX;
    endcase
    152: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    153: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd153;
      2: stateTransition = 11'd153;
      3: stateTransition = 11'd153;
      4: stateTransition = 11'd153;
      5: stateTransition = 11'd153;
      6: stateTransition = 11'd153;
      7: stateTransition = 11'd153;
      8: stateTransition = 11'd153;
      9: stateTransition = 11'd153;
      10: stateTransition = 11'd153;
      11: stateTransition = 11'd153;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd153;
      14: stateTransition = 11'd153;
      15: stateTransition = 11'd153;
      16: stateTransition = 11'd153;
      default: stateTransition = 11'bX;
    endcase
    154: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd154;
      2: stateTransition = 11'd154;
      3: stateTransition = 11'd154;
      4: stateTransition = 11'd154;
      5: stateTransition = 11'd154;
      6: stateTransition = 11'd154;
      7: stateTransition = 11'd154;
      8: stateTransition = 11'd154;
      9: stateTransition = 11'd154;
      10: stateTransition = 11'd154;
      11: stateTransition = 11'd154;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd154;
      14: stateTransition = 11'd154;
      15: stateTransition = 11'd154;
      16: stateTransition = 11'd154;
      default: stateTransition = 11'bX;
    endcase
    155: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd155;
      2: stateTransition = 11'd155;
      3: stateTransition = 11'd155;
      4: stateTransition = 11'd155;
      5: stateTransition = 11'd155;
      6: stateTransition = 11'd155;
      7: stateTransition = 11'd155;
      8: stateTransition = 11'd155;
      9: stateTransition = 11'd155;
      10: stateTransition = 11'd155;
      11: stateTransition = 11'd155;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd155;
      14: stateTransition = 11'd155;
      15: stateTransition = 11'd155;
      16: stateTransition = 11'd155;
      default: stateTransition = 11'bX;
    endcase
    156: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd156;
      2: stateTransition = 11'd156;
      3: stateTransition = 11'd156;
      4: stateTransition = 11'd156;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd156;
      7: stateTransition = 11'd156;
      8: stateTransition = 11'd156;
      9: stateTransition = 11'd156;
      10: stateTransition = 11'd156;
      11: stateTransition = 11'd156;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd156;
      14: stateTransition = 11'd156;
      15: stateTransition = 11'd156;
      16: stateTransition = 11'd156;
      default: stateTransition = 11'bX;
    endcase
    157: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd157;
      2: stateTransition = 11'd157;
      3: stateTransition = 11'd157;
      4: stateTransition = 11'd157;
      5: stateTransition = 11'd157;
      6: stateTransition = 11'd157;
      7: stateTransition = 11'd157;
      8: stateTransition = 11'd157;
      9: stateTransition = 11'd157;
      10: stateTransition = 11'd157;
      11: stateTransition = 11'd157;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd157;
      14: stateTransition = 11'd157;
      15: stateTransition = 11'd157;
      16: stateTransition = 11'd157;
      default: stateTransition = 11'bX;
    endcase
    158: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd158;
      2: stateTransition = 11'd158;
      3: stateTransition = 11'd158;
      4: stateTransition = 11'd158;
      5: stateTransition = 11'd158;
      6: stateTransition = 11'd158;
      7: stateTransition = 11'd158;
      8: stateTransition = 11'd158;
      9: stateTransition = 11'd158;
      10: stateTransition = 11'd158;
      11: stateTransition = 11'd158;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd158;
      14: stateTransition = 11'd158;
      15: stateTransition = 11'd158;
      16: stateTransition = 11'd158;
      default: stateTransition = 11'bX;
    endcase
    159: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd159;
      2: stateTransition = 11'd159;
      3: stateTransition = 11'd159;
      4: stateTransition = 11'd159;
      5: stateTransition = 11'd159;
      6: stateTransition = 11'd159;
      7: stateTransition = 11'd159;
      8: stateTransition = 11'd159;
      9: stateTransition = 11'd159;
      10: stateTransition = 11'd159;
      11: stateTransition = 11'd159;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd159;
      14: stateTransition = 11'd159;
      15: stateTransition = 11'd159;
      16: stateTransition = 11'd159;
      default: stateTransition = 11'bX;
    endcase
    160: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd160;
      2: stateTransition = 11'd160;
      3: stateTransition = 11'd160;
      4: stateTransition = 11'd160;
      5: stateTransition = 11'd160;
      6: stateTransition = 11'd160;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd160;
      9: stateTransition = 11'd160;
      10: stateTransition = 11'd160;
      11: stateTransition = 11'd160;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd160;
      14: stateTransition = 11'd160;
      15: stateTransition = 11'd160;
      16: stateTransition = 11'd160;
      default: stateTransition = 11'bX;
    endcase
    161: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd161;
      2: stateTransition = 11'd161;
      3: stateTransition = 11'd161;
      4: stateTransition = 11'd161;
      5: stateTransition = 11'd161;
      6: stateTransition = 11'd161;
      7: stateTransition = 11'd161;
      8: stateTransition = 11'd161;
      9: stateTransition = 11'd161;
      10: stateTransition = 11'd161;
      11: stateTransition = 11'd161;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd161;
      14: stateTransition = 11'd161;
      15: stateTransition = 11'd161;
      16: stateTransition = 11'd161;
      default: stateTransition = 11'bX;
    endcase
    162: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd162;
      2: stateTransition = 11'd162;
      3: stateTransition = 11'd162;
      4: stateTransition = 11'd162;
      5: stateTransition = 11'd162;
      6: stateTransition = 11'd162;
      7: stateTransition = 11'd162;
      8: stateTransition = 11'd162;
      9: stateTransition = 11'd162;
      10: stateTransition = 11'd162;
      11: stateTransition = 11'd162;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd162;
      14: stateTransition = 11'd162;
      15: stateTransition = 11'd162;
      16: stateTransition = 11'd162;
      default: stateTransition = 11'bX;
    endcase
    163: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd163;
      2: stateTransition = 11'd163;
      3: stateTransition = 11'd163;
      4: stateTransition = 11'd163;
      5: stateTransition = 11'd163;
      6: stateTransition = 11'd163;
      7: stateTransition = 11'd163;
      8: stateTransition = 11'd163;
      9: stateTransition = 11'd163;
      10: stateTransition = 11'd163;
      11: stateTransition = 11'd163;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd163;
      14: stateTransition = 11'd163;
      15: stateTransition = 11'd163;
      16: stateTransition = 11'd163;
      default: stateTransition = 11'bX;
    endcase
    164: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd164;
      2: stateTransition = 11'd164;
      3: stateTransition = 11'd164;
      4: stateTransition = 11'd164;
      5: stateTransition = 11'd164;
      6: stateTransition = 11'd164;
      7: stateTransition = 11'd164;
      8: stateTransition = 11'd164;
      9: stateTransition = 11'd164;
      10: stateTransition = 11'd164;
      11: stateTransition = 11'd164;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd164;
      14: stateTransition = 11'd164;
      15: stateTransition = 11'd164;
      16: stateTransition = 11'd164;
      default: stateTransition = 11'bX;
    endcase
    165: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd165;
      2: stateTransition = 11'd165;
      3: stateTransition = 11'd165;
      4: stateTransition = 11'd165;
      5: stateTransition = 11'd165;
      6: stateTransition = 11'd165;
      7: stateTransition = 11'd165;
      8: stateTransition = 11'd165;
      9: stateTransition = 11'd165;
      10: stateTransition = 11'd165;
      11: stateTransition = 11'd165;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd165;
      14: stateTransition = 11'd165;
      15: stateTransition = 11'd165;
      16: stateTransition = 11'd165;
      default: stateTransition = 11'bX;
    endcase
    166: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd166;
      2: stateTransition = 11'd166;
      3: stateTransition = 11'd166;
      4: stateTransition = 11'd166;
      5: stateTransition = 11'd166;
      6: stateTransition = 11'd166;
      7: stateTransition = 11'd166;
      8: stateTransition = 11'd166;
      9: stateTransition = 11'd166;
      10: stateTransition = 11'd166;
      11: stateTransition = 11'd166;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd166;
      14: stateTransition = 11'd166;
      15: stateTransition = 11'd166;
      16: stateTransition = 11'd166;
      default: stateTransition = 11'bX;
    endcase
    167: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd167;
      2: stateTransition = 11'd167;
      3: stateTransition = 11'd167;
      4: stateTransition = 11'd167;
      5: stateTransition = 11'd167;
      6: stateTransition = 11'd167;
      7: stateTransition = 11'd167;
      8: stateTransition = 11'd167;
      9: stateTransition = 11'd167;
      10: stateTransition = 11'd167;
      11: stateTransition = 11'd167;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd167;
      14: stateTransition = 11'd167;
      15: stateTransition = 11'd167;
      16: stateTransition = 11'd167;
      default: stateTransition = 11'bX;
    endcase
    168: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd168;
      2: stateTransition = 11'd168;
      3: stateTransition = 11'd168;
      4: stateTransition = 11'd168;
      5: stateTransition = 11'd168;
      6: stateTransition = 11'd168;
      7: stateTransition = 11'd168;
      8: stateTransition = 11'd168;
      9: stateTransition = 11'd168;
      10: stateTransition = 11'd168;
      11: stateTransition = 11'd168;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd168;
      14: stateTransition = 11'd168;
      15: stateTransition = 11'd168;
      16: stateTransition = 11'd168;
      default: stateTransition = 11'bX;
    endcase
    169: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd169;
      2: stateTransition = 11'd169;
      3: stateTransition = 11'd169;
      4: stateTransition = 11'd169;
      5: stateTransition = 11'd169;
      6: stateTransition = 11'd169;
      7: stateTransition = 11'd169;
      8: stateTransition = 11'd169;
      9: stateTransition = 11'd169;
      10: stateTransition = 11'd169;
      11: stateTransition = 11'd169;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd169;
      14: stateTransition = 11'd169;
      15: stateTransition = 11'd169;
      16: stateTransition = 11'd169;
      default: stateTransition = 11'bX;
    endcase
    170: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd170;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd170;
      5: stateTransition = 11'd170;
      6: stateTransition = 11'd170;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd170;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    171: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd171;
      2: stateTransition = 11'd171;
      3: stateTransition = 11'd171;
      4: stateTransition = 11'd171;
      5: stateTransition = 11'd171;
      6: stateTransition = 11'd171;
      7: stateTransition = 11'd171;
      8: stateTransition = 11'd171;
      9: stateTransition = 11'd171;
      10: stateTransition = 11'd171;
      11: stateTransition = 11'd171;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd171;
      14: stateTransition = 11'd171;
      15: stateTransition = 11'd171;
      16: stateTransition = 11'd171;
      default: stateTransition = 11'bX;
    endcase
    172: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd172;
      5: stateTransition = 11'd172;
      6: stateTransition = 11'd172;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd172;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    173: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd173;
      2: stateTransition = 11'd173;
      3: stateTransition = 11'd173;
      4: stateTransition = 11'd173;
      5: stateTransition = 11'd173;
      6: stateTransition = 11'd173;
      7: stateTransition = 11'd173;
      8: stateTransition = 11'd173;
      9: stateTransition = 11'd173;
      10: stateTransition = 11'd173;
      11: stateTransition = 11'd173;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd173;
      14: stateTransition = 11'd173;
      15: stateTransition = 11'd173;
      16: stateTransition = 11'd173;
      default: stateTransition = 11'bX;
    endcase
    174: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd174;
      2: stateTransition = 11'd174;
      3: stateTransition = 11'd174;
      4: stateTransition = 11'd174;
      5: stateTransition = 11'd174;
      6: stateTransition = 11'd174;
      7: stateTransition = 11'd174;
      8: stateTransition = 11'd174;
      9: stateTransition = 11'd174;
      10: stateTransition = 11'd174;
      11: stateTransition = 11'd174;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd174;
      14: stateTransition = 11'd174;
      15: stateTransition = 11'd174;
      16: stateTransition = 11'd174;
      default: stateTransition = 11'bX;
    endcase
    175: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd175;
      2: stateTransition = 11'd175;
      3: stateTransition = 11'd175;
      4: stateTransition = 11'd175;
      5: stateTransition = 11'd175;
      6: stateTransition = 11'd175;
      7: stateTransition = 11'd175;
      8: stateTransition = 11'd175;
      9: stateTransition = 11'd175;
      10: stateTransition = 11'd175;
      11: stateTransition = 11'd175;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd175;
      14: stateTransition = 11'd175;
      15: stateTransition = 11'd175;
      16: stateTransition = 11'd175;
      default: stateTransition = 11'bX;
    endcase
    176: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd176;
      2: stateTransition = 11'd176;
      3: stateTransition = 11'd176;
      4: stateTransition = 11'd176;
      5: stateTransition = 11'd176;
      6: stateTransition = 11'd176;
      7: stateTransition = 11'd176;
      8: stateTransition = 11'd176;
      9: stateTransition = 11'd176;
      10: stateTransition = 11'd176;
      11: stateTransition = 11'd176;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd176;
      14: stateTransition = 11'd176;
      15: stateTransition = 11'd176;
      16: stateTransition = 11'd176;
      default: stateTransition = 11'bX;
    endcase
    177: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd177;
      2: stateTransition = 11'd177;
      3: stateTransition = 11'd177;
      4: stateTransition = 11'd177;
      5: stateTransition = 11'd177;
      6: stateTransition = 11'd177;
      7: stateTransition = 11'd177;
      8: stateTransition = 11'd177;
      9: stateTransition = 11'd177;
      10: stateTransition = 11'd177;
      11: stateTransition = 11'd177;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd177;
      14: stateTransition = 11'd177;
      15: stateTransition = 11'd177;
      16: stateTransition = 11'd177;
      default: stateTransition = 11'bX;
    endcase
    178: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd178;
      2: stateTransition = 11'd178;
      3: stateTransition = 11'd178;
      4: stateTransition = 11'd178;
      5: stateTransition = 11'd178;
      6: stateTransition = 11'd178;
      7: stateTransition = 11'd178;
      8: stateTransition = 11'd178;
      9: stateTransition = 11'd178;
      10: stateTransition = 11'd178;
      11: stateTransition = 11'd178;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd178;
      14: stateTransition = 11'd178;
      15: stateTransition = 11'd178;
      16: stateTransition = 11'd178;
      default: stateTransition = 11'bX;
    endcase
    179: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd179;
      2: stateTransition = 11'd179;
      3: stateTransition = 11'd179;
      4: stateTransition = 11'd179;
      5: stateTransition = 11'd179;
      6: stateTransition = 11'd179;
      7: stateTransition = 11'd179;
      8: stateTransition = 11'd179;
      9: stateTransition = 11'd179;
      10: stateTransition = 11'd179;
      11: stateTransition = 11'd179;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd179;
      14: stateTransition = 11'd179;
      15: stateTransition = 11'd179;
      16: stateTransition = 11'd179;
      default: stateTransition = 11'bX;
    endcase
    180: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd180;
      2: stateTransition = 11'd180;
      3: stateTransition = 11'd180;
      4: stateTransition = 11'd180;
      5: stateTransition = 11'd180;
      6: stateTransition = 11'd180;
      7: stateTransition = 11'd180;
      8: stateTransition = 11'd180;
      9: stateTransition = 11'd180;
      10: stateTransition = 11'd180;
      11: stateTransition = 11'd180;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd180;
      14: stateTransition = 11'd180;
      15: stateTransition = 11'd180;
      16: stateTransition = 11'd180;
      default: stateTransition = 11'bX;
    endcase
    181: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd181;
      2: stateTransition = 11'd181;
      3: stateTransition = 11'd181;
      4: stateTransition = 11'd181;
      5: stateTransition = 11'd181;
      6: stateTransition = 11'd181;
      7: stateTransition = 11'd181;
      8: stateTransition = 11'd181;
      9: stateTransition = 11'd181;
      10: stateTransition = 11'd181;
      11: stateTransition = 11'd181;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd181;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd181;
      16: stateTransition = 11'd181;
      default: stateTransition = 11'bX;
    endcase
    182: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd182;
      2: stateTransition = 11'd182;
      3: stateTransition = 11'd182;
      4: stateTransition = 11'd182;
      5: stateTransition = 11'd182;
      6: stateTransition = 11'd182;
      7: stateTransition = 11'd182;
      8: stateTransition = 11'd182;
      9: stateTransition = 11'd182;
      10: stateTransition = 11'd182;
      11: stateTransition = 11'd182;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd182;
      14: stateTransition = 11'd182;
      15: stateTransition = 11'd182;
      16: stateTransition = 11'd182;
      default: stateTransition = 11'bX;
    endcase
    183: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd183;
      2: stateTransition = 11'd183;
      3: stateTransition = 11'd183;
      4: stateTransition = 11'd183;
      5: stateTransition = 11'd183;
      6: stateTransition = 11'd183;
      7: stateTransition = 11'd183;
      8: stateTransition = 11'd183;
      9: stateTransition = 11'd183;
      10: stateTransition = 11'd183;
      11: stateTransition = 11'd183;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd183;
      14: stateTransition = 11'd183;
      15: stateTransition = 11'd183;
      16: stateTransition = 11'd183;
      default: stateTransition = 11'bX;
    endcase
    184: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd184;
      2: stateTransition = 11'd184;
      3: stateTransition = 11'd184;
      4: stateTransition = 11'd184;
      5: stateTransition = 11'd184;
      6: stateTransition = 11'd184;
      7: stateTransition = 11'd184;
      8: stateTransition = 11'd184;
      9: stateTransition = 11'd184;
      10: stateTransition = 11'd184;
      11: stateTransition = 11'd184;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd184;
      14: stateTransition = 11'd184;
      15: stateTransition = 11'd184;
      16: stateTransition = 11'd184;
      default: stateTransition = 11'bX;
    endcase
    185: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd185;
      2: stateTransition = 11'd185;
      3: stateTransition = 11'd185;
      4: stateTransition = 11'd185;
      5: stateTransition = 11'd185;
      6: stateTransition = 11'd185;
      7: stateTransition = 11'd185;
      8: stateTransition = 11'd185;
      9: stateTransition = 11'd185;
      10: stateTransition = 11'd185;
      11: stateTransition = 11'd185;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd185;
      14: stateTransition = 11'd185;
      15: stateTransition = 11'd185;
      16: stateTransition = 11'd185;
      default: stateTransition = 11'bX;
    endcase
    186: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    187: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd187;
      2: stateTransition = 11'd187;
      3: stateTransition = 11'd187;
      4: stateTransition = 11'd187;
      5: stateTransition = 11'd187;
      6: stateTransition = 11'd187;
      7: stateTransition = 11'd187;
      8: stateTransition = 11'd187;
      9: stateTransition = 11'd187;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd187;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd187;
      14: stateTransition = 11'd187;
      15: stateTransition = 11'd187;
      16: stateTransition = 11'd187;
      default: stateTransition = 11'bX;
    endcase
    188: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd188;
      2: stateTransition = 11'd188;
      3: stateTransition = 11'd188;
      4: stateTransition = 11'd188;
      5: stateTransition = 11'd188;
      6: stateTransition = 11'd188;
      7: stateTransition = 11'd188;
      8: stateTransition = 11'd188;
      9: stateTransition = 11'd188;
      10: stateTransition = 11'd188;
      11: stateTransition = 11'd188;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd188;
      14: stateTransition = 11'd188;
      15: stateTransition = 11'd188;
      16: stateTransition = 11'd188;
      default: stateTransition = 11'bX;
    endcase
    189: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd189;
      2: stateTransition = 11'd189;
      3: stateTransition = 11'd189;
      4: stateTransition = 11'd189;
      5: stateTransition = 11'd189;
      6: stateTransition = 11'd189;
      7: stateTransition = 11'd189;
      8: stateTransition = 11'd189;
      9: stateTransition = 11'd189;
      10: stateTransition = 11'd189;
      11: stateTransition = 11'd189;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd189;
      14: stateTransition = 11'd189;
      15: stateTransition = 11'd189;
      16: stateTransition = 11'd189;
      default: stateTransition = 11'bX;
    endcase
    190: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd190;
      2: stateTransition = 11'd190;
      3: stateTransition = 11'd190;
      4: stateTransition = 11'd190;
      5: stateTransition = 11'd190;
      6: stateTransition = 11'd190;
      7: stateTransition = 11'd190;
      8: stateTransition = 11'd190;
      9: stateTransition = 11'd190;
      10: stateTransition = 11'd190;
      11: stateTransition = 11'd190;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd190;
      14: stateTransition = 11'd190;
      15: stateTransition = 11'd190;
      16: stateTransition = 11'd190;
      default: stateTransition = 11'bX;
    endcase
    191: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd191;
      2: stateTransition = 11'd191;
      3: stateTransition = 11'd191;
      4: stateTransition = 11'd191;
      5: stateTransition = 11'd191;
      6: stateTransition = 11'd191;
      7: stateTransition = 11'd191;
      8: stateTransition = 11'd191;
      9: stateTransition = 11'd191;
      10: stateTransition = 11'd191;
      11: stateTransition = 11'd191;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd191;
      14: stateTransition = 11'd191;
      15: stateTransition = 11'd191;
      16: stateTransition = 11'd191;
      default: stateTransition = 11'bX;
    endcase
    192: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd192;
      2: stateTransition = 11'd192;
      3: stateTransition = 11'd192;
      4: stateTransition = 11'd192;
      5: stateTransition = 11'd192;
      6: stateTransition = 11'd192;
      7: stateTransition = 11'd192;
      8: stateTransition = 11'd192;
      9: stateTransition = 11'd192;
      10: stateTransition = 11'd192;
      11: stateTransition = 11'd192;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd192;
      14: stateTransition = 11'd192;
      15: stateTransition = 11'd192;
      16: stateTransition = 11'd192;
      default: stateTransition = 11'bX;
    endcase
    193: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd193;
      2: stateTransition = 11'd193;
      3: stateTransition = 11'd193;
      4: stateTransition = 11'd193;
      5: stateTransition = 11'd193;
      6: stateTransition = 11'd193;
      7: stateTransition = 11'd193;
      8: stateTransition = 11'd193;
      9: stateTransition = 11'd193;
      10: stateTransition = 11'd193;
      11: stateTransition = 11'd193;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd193;
      14: stateTransition = 11'd193;
      15: stateTransition = 11'd193;
      16: stateTransition = 11'd193;
      default: stateTransition = 11'bX;
    endcase
    194: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd194;
      2: stateTransition = 11'd194;
      3: stateTransition = 11'd194;
      4: stateTransition = 11'd194;
      5: stateTransition = 11'd194;
      6: stateTransition = 11'd194;
      7: stateTransition = 11'd194;
      8: stateTransition = 11'd194;
      9: stateTransition = 11'd194;
      10: stateTransition = 11'd194;
      11: stateTransition = 11'd194;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd194;
      14: stateTransition = 11'd194;
      15: stateTransition = 11'd194;
      16: stateTransition = 11'd194;
      default: stateTransition = 11'bX;
    endcase
    195: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd195;
      3: stateTransition = 11'd195;
      4: stateTransition = 11'd195;
      5: stateTransition = 11'd195;
      6: stateTransition = 11'd195;
      7: stateTransition = 11'd195;
      8: stateTransition = 11'd195;
      9: stateTransition = 11'd195;
      10: stateTransition = 11'd195;
      11: stateTransition = 11'd195;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd195;
      14: stateTransition = 11'd195;
      15: stateTransition = 11'd195;
      16: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    196: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd196;
      2: stateTransition = 11'd196;
      3: stateTransition = 11'd196;
      4: stateTransition = 11'd196;
      5: stateTransition = 11'd196;
      6: stateTransition = 11'd196;
      7: stateTransition = 11'd196;
      8: stateTransition = 11'd196;
      9: stateTransition = 11'd196;
      10: stateTransition = 11'd196;
      11: stateTransition = 11'd196;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd196;
      14: stateTransition = 11'd196;
      15: stateTransition = 11'd196;
      16: stateTransition = 11'd196;
      default: stateTransition = 11'bX;
    endcase
    197: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd197;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd197;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd197;
      8: stateTransition = 11'd197;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      default: stateTransition = 11'bX;
    endcase
    198: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd198;
      2: stateTransition = 11'd198;
      3: stateTransition = 11'd198;
      4: stateTransition = 11'd198;
      5: stateTransition = 11'd198;
      6: stateTransition = 11'd198;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd198;
      10: stateTransition = 11'd198;
      11: stateTransition = 11'd198;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd198;
      14: stateTransition = 11'd198;
      15: stateTransition = 11'd198;
      16: stateTransition = 11'd198;
      default: stateTransition = 11'bX;
    endcase
    199: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd199;
      2: stateTransition = 11'd199;
      3: stateTransition = 11'd199;
      4: stateTransition = 11'd199;
      5: stateTransition = 11'd199;
      6: stateTransition = 11'd199;
      7: stateTransition = 11'd199;
      8: stateTransition = 11'd199;
      9: stateTransition = 11'd199;
      10: stateTransition = 11'd199;
      11: stateTransition = 11'd199;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd199;
      14: stateTransition = 11'd199;
      15: stateTransition = 11'd199;
      16: stateTransition = 11'd199;
      default: stateTransition = 11'bX;
    endcase
    200: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd200;
      2: stateTransition = 11'd200;
      3: stateTransition = 11'd200;
      4: stateTransition = 11'd200;
      5: stateTransition = 11'd200;
      6: stateTransition = 11'd200;
      7: stateTransition = 11'd200;
      8: stateTransition = 11'd200;
      9: stateTransition = 11'd200;
      10: stateTransition = 11'd200;
      11: stateTransition = 11'd200;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd200;
      14: stateTransition = 11'd200;
      15: stateTransition = 11'd200;
      16: stateTransition = 11'd200;
      default: stateTransition = 11'bX;
    endcase
    201: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd201;
      2: stateTransition = 11'd201;
      3: stateTransition = 11'd201;
      4: stateTransition = 11'd201;
      5: stateTransition = 11'd201;
      6: stateTransition = 11'd201;
      7: stateTransition = 11'd201;
      8: stateTransition = 11'd201;
      9: stateTransition = 11'd201;
      10: stateTransition = 11'd201;
      11: stateTransition = 11'd201;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd201;
      14: stateTransition = 11'd201;
      15: stateTransition = 11'd201;
      16: stateTransition = 11'd201;
      default: stateTransition = 11'bX;
    endcase
    202: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd202;
      2: stateTransition = 11'd202;
      3: stateTransition = 11'd202;
      4: stateTransition = 11'd202;
      5: stateTransition = 11'd202;
      6: stateTransition = 11'd202;
      7: stateTransition = 11'd202;
      8: stateTransition = 11'd202;
      9: stateTransition = 11'd202;
      10: stateTransition = 11'd202;
      11: stateTransition = 11'd202;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd202;
      14: stateTransition = 11'd202;
      15: stateTransition = 11'd202;
      16: stateTransition = 11'd202;
      default: stateTransition = 11'bX;
    endcase
    203: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd203;
      2: stateTransition = 11'd203;
      3: stateTransition = 11'd203;
      4: stateTransition = 11'd203;
      5: stateTransition = 11'd203;
      6: stateTransition = 11'd203;
      7: stateTransition = 11'd203;
      8: stateTransition = 11'd203;
      9: stateTransition = 11'd203;
      10: stateTransition = 11'd203;
      11: stateTransition = 11'd203;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd203;
      14: stateTransition = 11'd203;
      15: stateTransition = 11'd203;
      16: stateTransition = 11'd203;
      default: stateTransition = 11'bX;
    endcase
    204: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd204;
      2: stateTransition = 11'd204;
      3: stateTransition = 11'd204;
      4: stateTransition = 11'd204;
      5: stateTransition = 11'd204;
      6: stateTransition = 11'd204;
      7: stateTransition = 11'd204;
      8: stateTransition = 11'd204;
      9: stateTransition = 11'd204;
      10: stateTransition = 11'd204;
      11: stateTransition = 11'd204;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd204;
      14: stateTransition = 11'd204;
      15: stateTransition = 11'd204;
      16: stateTransition = 11'd204;
      default: stateTransition = 11'bX;
    endcase
    205: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd205;
      2: stateTransition = 11'd205;
      3: stateTransition = 11'd205;
      4: stateTransition = 11'd205;
      5: stateTransition = 11'd205;
      6: stateTransition = 11'd205;
      7: stateTransition = 11'd205;
      8: stateTransition = 11'd205;
      9: stateTransition = 11'd205;
      10: stateTransition = 11'd205;
      11: stateTransition = 11'd205;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd205;
      14: stateTransition = 11'd205;
      15: stateTransition = 11'd205;
      16: stateTransition = 11'd205;
      default: stateTransition = 11'bX;
    endcase
    206: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd206;
      2: stateTransition = 11'd206;
      3: stateTransition = 11'd206;
      4: stateTransition = 11'd206;
      5: stateTransition = 11'd206;
      6: stateTransition = 11'd206;
      7: stateTransition = 11'd206;
      8: stateTransition = 11'd206;
      9: stateTransition = 11'd206;
      10: stateTransition = 11'd206;
      11: stateTransition = 11'd206;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd206;
      14: stateTransition = 11'd206;
      15: stateTransition = 11'd206;
      16: stateTransition = 11'd206;
      default: stateTransition = 11'bX;
    endcase
    207: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd207;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd207;
      5: stateTransition = 11'd207;
      6: stateTransition = 11'd207;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd207;
      9: stateTransition = 11'd207;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd207;
      14: stateTransition = 11'd207;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    208: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd208;
      2: stateTransition = 11'd208;
      3: stateTransition = 11'd208;
      4: stateTransition = 11'd208;
      5: stateTransition = 11'd208;
      6: stateTransition = 11'd208;
      7: stateTransition = 11'd208;
      8: stateTransition = 11'd208;
      9: stateTransition = 11'd208;
      10: stateTransition = 11'd208;
      11: stateTransition = 11'd208;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd208;
      14: stateTransition = 11'd208;
      15: stateTransition = 11'd208;
      16: stateTransition = 11'd208;
      default: stateTransition = 11'bX;
    endcase
    209: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd209;
      2: stateTransition = 11'd209;
      3: stateTransition = 11'd209;
      4: stateTransition = 11'd209;
      5: stateTransition = 11'd209;
      6: stateTransition = 11'd209;
      7: stateTransition = 11'd209;
      8: stateTransition = 11'd209;
      9: stateTransition = 11'd209;
      10: stateTransition = 11'd209;
      11: stateTransition = 11'd209;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd209;
      14: stateTransition = 11'd209;
      15: stateTransition = 11'd209;
      16: stateTransition = 11'd209;
      default: stateTransition = 11'bX;
    endcase
    210: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd210;
      2: stateTransition = 11'd210;
      3: stateTransition = 11'd210;
      4: stateTransition = 11'd210;
      5: stateTransition = 11'd210;
      6: stateTransition = 11'd210;
      7: stateTransition = 11'd210;
      8: stateTransition = 11'd210;
      9: stateTransition = 11'd210;
      10: stateTransition = 11'd210;
      11: stateTransition = 11'd210;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd210;
      14: stateTransition = 11'd210;
      15: stateTransition = 11'd210;
      16: stateTransition = 11'd210;
      default: stateTransition = 11'bX;
    endcase
    211: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd211;
      2: stateTransition = 11'd211;
      3: stateTransition = 11'd211;
      4: stateTransition = 11'd211;
      5: stateTransition = 11'd211;
      6: stateTransition = 11'd211;
      7: stateTransition = 11'd211;
      8: stateTransition = 11'd211;
      9: stateTransition = 11'd211;
      10: stateTransition = 11'd211;
      11: stateTransition = 11'd211;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd211;
      14: stateTransition = 11'd211;
      15: stateTransition = 11'd211;
      16: stateTransition = 11'd211;
      default: stateTransition = 11'bX;
    endcase
    212: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd212;
      2: stateTransition = 11'd212;
      3: stateTransition = 11'd212;
      4: stateTransition = 11'd212;
      5: stateTransition = 11'd212;
      6: stateTransition = 11'd212;
      7: stateTransition = 11'd212;
      8: stateTransition = 11'd212;
      9: stateTransition = 11'd212;
      10: stateTransition = 11'd212;
      11: stateTransition = 11'd212;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd212;
      14: stateTransition = 11'd212;
      15: stateTransition = 11'd212;
      16: stateTransition = 11'd212;
      default: stateTransition = 11'bX;
    endcase
    213: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd213;
      2: stateTransition = 11'd213;
      3: stateTransition = 11'd213;
      4: stateTransition = 11'd213;
      5: stateTransition = 11'd213;
      6: stateTransition = 11'd213;
      7: stateTransition = 11'd213;
      8: stateTransition = 11'd213;
      9: stateTransition = 11'd213;
      10: stateTransition = 11'd213;
      11: stateTransition = 11'd213;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd213;
      14: stateTransition = 11'd213;
      15: stateTransition = 11'd213;
      16: stateTransition = 11'd213;
      default: stateTransition = 11'bX;
    endcase
    214: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd214;
      2: stateTransition = 11'd214;
      3: stateTransition = 11'd214;
      4: stateTransition = 11'd214;
      5: stateTransition = 11'd214;
      6: stateTransition = 11'd214;
      7: stateTransition = 11'd214;
      8: stateTransition = 11'd214;
      9: stateTransition = 11'd214;
      10: stateTransition = 11'd214;
      11: stateTransition = 11'd214;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd214;
      14: stateTransition = 11'd214;
      15: stateTransition = 11'd214;
      16: stateTransition = 11'd214;
      default: stateTransition = 11'bX;
    endcase
    215: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd215;
      2: stateTransition = 11'd215;
      3: stateTransition = 11'd215;
      4: stateTransition = 11'd215;
      5: stateTransition = 11'd215;
      6: stateTransition = 11'd215;
      7: stateTransition = 11'd215;
      8: stateTransition = 11'd215;
      9: stateTransition = 11'd215;
      10: stateTransition = 11'd215;
      11: stateTransition = 11'd215;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd215;
      14: stateTransition = 11'd215;
      15: stateTransition = 11'd215;
      16: stateTransition = 11'd215;
      default: stateTransition = 11'bX;
    endcase
    216: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd216;
      2: stateTransition = 11'd216;
      3: stateTransition = 11'd216;
      4: stateTransition = 11'd216;
      5: stateTransition = 11'd216;
      6: stateTransition = 11'd216;
      7: stateTransition = 11'd216;
      8: stateTransition = 11'd216;
      9: stateTransition = 11'd216;
      10: stateTransition = 11'd216;
      11: stateTransition = 11'd216;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd216;
      14: stateTransition = 11'd216;
      15: stateTransition = 11'd216;
      16: stateTransition = 11'd216;
      default: stateTransition = 11'bX;
    endcase
    217: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd217;
      2: stateTransition = 11'd217;
      3: stateTransition = 11'd217;
      4: stateTransition = 11'd217;
      5: stateTransition = 11'd217;
      6: stateTransition = 11'd217;
      7: stateTransition = 11'd217;
      8: stateTransition = 11'd217;
      9: stateTransition = 11'd217;
      10: stateTransition = 11'd217;
      11: stateTransition = 11'd217;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd217;
      14: stateTransition = 11'd217;
      15: stateTransition = 11'd217;
      16: stateTransition = 11'd217;
      default: stateTransition = 11'bX;
    endcase
    218: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd218;
      2: stateTransition = 11'd218;
      3: stateTransition = 11'd218;
      4: stateTransition = 11'd218;
      5: stateTransition = 11'd218;
      6: stateTransition = 11'd218;
      7: stateTransition = 11'd218;
      8: stateTransition = 11'd218;
      9: stateTransition = 11'd218;
      10: stateTransition = 11'd218;
      11: stateTransition = 11'd218;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd218;
      14: stateTransition = 11'd218;
      15: stateTransition = 11'd218;
      16: stateTransition = 11'd218;
      default: stateTransition = 11'bX;
    endcase
    219: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd219;
      2: stateTransition = 11'd219;
      3: stateTransition = 11'd219;
      4: stateTransition = 11'd219;
      5: stateTransition = 11'd219;
      6: stateTransition = 11'd219;
      7: stateTransition = 11'd219;
      8: stateTransition = 11'd219;
      9: stateTransition = 11'd219;
      10: stateTransition = 11'd219;
      11: stateTransition = 11'd219;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd219;
      14: stateTransition = 11'd219;
      15: stateTransition = 11'd219;
      16: stateTransition = 11'd219;
      default: stateTransition = 11'bX;
    endcase
    220: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd220;
      2: stateTransition = 11'd220;
      3: stateTransition = 11'd220;
      4: stateTransition = 11'd220;
      5: stateTransition = 11'd220;
      6: stateTransition = 11'd220;
      7: stateTransition = 11'd220;
      8: stateTransition = 11'd220;
      9: stateTransition = 11'd220;
      10: stateTransition = 11'd220;
      11: stateTransition = 11'd220;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd220;
      14: stateTransition = 11'd220;
      15: stateTransition = 11'd220;
      16: stateTransition = 11'd220;
      default: stateTransition = 11'bX;
    endcase
    221: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd221;
      2: stateTransition = 11'd221;
      3: stateTransition = 11'd221;
      4: stateTransition = 11'd221;
      5: stateTransition = 11'd221;
      6: stateTransition = 11'd221;
      7: stateTransition = 11'd221;
      8: stateTransition = 11'd221;
      9: stateTransition = 11'd221;
      10: stateTransition = 11'd221;
      11: stateTransition = 11'd221;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd221;
      14: stateTransition = 11'd221;
      15: stateTransition = 11'd221;
      16: stateTransition = 11'd221;
      default: stateTransition = 11'bX;
    endcase
    222: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd222;
      2: stateTransition = 11'd222;
      3: stateTransition = 11'd222;
      4: stateTransition = 11'd222;
      5: stateTransition = 11'd222;
      6: stateTransition = 11'd222;
      7: stateTransition = 11'd222;
      8: stateTransition = 11'd222;
      9: stateTransition = 11'd222;
      10: stateTransition = 11'd222;
      11: stateTransition = 11'd222;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd222;
      14: stateTransition = 11'd222;
      15: stateTransition = 11'd222;
      16: stateTransition = 11'd222;
      default: stateTransition = 11'bX;
    endcase
    223: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd223;
      2: stateTransition = 11'd223;
      3: stateTransition = 11'd223;
      4: stateTransition = 11'd223;
      5: stateTransition = 11'd223;
      6: stateTransition = 11'd223;
      7: stateTransition = 11'd223;
      8: stateTransition = 11'd223;
      9: stateTransition = 11'd223;
      10: stateTransition = 11'd223;
      11: stateTransition = 11'd223;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd223;
      14: stateTransition = 11'd223;
      15: stateTransition = 11'd223;
      16: stateTransition = 11'd223;
      default: stateTransition = 11'bX;
    endcase
    224: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd224;
      2: stateTransition = 11'd224;
      3: stateTransition = 11'd224;
      4: stateTransition = 11'd224;
      5: stateTransition = 11'd224;
      6: stateTransition = 11'd224;
      7: stateTransition = 11'd224;
      8: stateTransition = 11'd224;
      9: stateTransition = 11'd224;
      10: stateTransition = 11'd224;
      11: stateTransition = 11'd224;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd224;
      14: stateTransition = 11'd224;
      15: stateTransition = 11'd224;
      16: stateTransition = 11'd224;
      default: stateTransition = 11'bX;
    endcase
    225: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd225;
      2: stateTransition = 11'd225;
      3: stateTransition = 11'd225;
      4: stateTransition = 11'd225;
      5: stateTransition = 11'd225;
      6: stateTransition = 11'd225;
      7: stateTransition = 11'd225;
      8: stateTransition = 11'd225;
      9: stateTransition = 11'd225;
      10: stateTransition = 11'd225;
      11: stateTransition = 11'd225;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd225;
      14: stateTransition = 11'd225;
      15: stateTransition = 11'd225;
      16: stateTransition = 11'd225;
      default: stateTransition = 11'bX;
    endcase
    226: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd226;
      2: stateTransition = 11'd226;
      3: stateTransition = 11'd226;
      4: stateTransition = 11'd226;
      5: stateTransition = 11'd226;
      6: stateTransition = 11'd226;
      7: stateTransition = 11'd226;
      8: stateTransition = 11'd226;
      9: stateTransition = 11'd226;
      10: stateTransition = 11'd226;
      11: stateTransition = 11'd226;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd226;
      14: stateTransition = 11'd226;
      15: stateTransition = 11'd226;
      16: stateTransition = 11'd226;
      default: stateTransition = 11'bX;
    endcase
    227: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd227;
      2: stateTransition = 11'd227;
      3: stateTransition = 11'd227;
      4: stateTransition = 11'd227;
      5: stateTransition = 11'd227;
      6: stateTransition = 11'd227;
      7: stateTransition = 11'd227;
      8: stateTransition = 11'd227;
      9: stateTransition = 11'd227;
      10: stateTransition = 11'd227;
      11: stateTransition = 11'd227;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd227;
      14: stateTransition = 11'd227;
      15: stateTransition = 11'd227;
      16: stateTransition = 11'd227;
      default: stateTransition = 11'bX;
    endcase
    228: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd228;
      2: stateTransition = 11'd228;
      3: stateTransition = 11'd228;
      4: stateTransition = 11'd228;
      5: stateTransition = 11'd228;
      6: stateTransition = 11'd228;
      7: stateTransition = 11'd228;
      8: stateTransition = 11'd228;
      9: stateTransition = 11'd228;
      10: stateTransition = 11'd228;
      11: stateTransition = 11'd228;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd228;
      14: stateTransition = 11'd228;
      15: stateTransition = 11'd228;
      16: stateTransition = 11'd228;
      default: stateTransition = 11'bX;
    endcase
    229: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd229;
      2: stateTransition = 11'd229;
      3: stateTransition = 11'd229;
      4: stateTransition = 11'd229;
      5: stateTransition = 11'd229;
      6: stateTransition = 11'd229;
      7: stateTransition = 11'd229;
      8: stateTransition = 11'd229;
      9: stateTransition = 11'd229;
      10: stateTransition = 11'd229;
      11: stateTransition = 11'd229;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd229;
      14: stateTransition = 11'd229;
      15: stateTransition = 11'd229;
      16: stateTransition = 11'd229;
      default: stateTransition = 11'bX;
    endcase
    230: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd230;
      2: stateTransition = 11'd230;
      3: stateTransition = 11'd230;
      4: stateTransition = 11'd230;
      5: stateTransition = 11'd230;
      6: stateTransition = 11'd230;
      7: stateTransition = 11'd230;
      8: stateTransition = 11'd230;
      9: stateTransition = 11'd230;
      10: stateTransition = 11'd230;
      11: stateTransition = 11'd230;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd230;
      14: stateTransition = 11'd230;
      15: stateTransition = 11'd230;
      16: stateTransition = 11'd230;
      default: stateTransition = 11'bX;
    endcase
    231: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd231;
      2: stateTransition = 11'd231;
      3: stateTransition = 11'd231;
      4: stateTransition = 11'd231;
      5: stateTransition = 11'd231;
      6: stateTransition = 11'd231;
      7: stateTransition = 11'd231;
      8: stateTransition = 11'd231;
      9: stateTransition = 11'd231;
      10: stateTransition = 11'd231;
      11: stateTransition = 11'd231;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd231;
      14: stateTransition = 11'd231;
      15: stateTransition = 11'd231;
      16: stateTransition = 11'd231;
      default: stateTransition = 11'bX;
    endcase
    232: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd232;
      2: stateTransition = 11'd232;
      3: stateTransition = 11'd232;
      4: stateTransition = 11'd232;
      5: stateTransition = 11'd232;
      6: stateTransition = 11'd232;
      7: stateTransition = 11'd232;
      8: stateTransition = 11'd232;
      9: stateTransition = 11'd232;
      10: stateTransition = 11'd232;
      11: stateTransition = 11'd232;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd232;
      14: stateTransition = 11'd232;
      15: stateTransition = 11'd232;
      16: stateTransition = 11'd232;
      default: stateTransition = 11'bX;
    endcase
    233: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd233;
      2: stateTransition = 11'd233;
      3: stateTransition = 11'd233;
      4: stateTransition = 11'd233;
      5: stateTransition = 11'd233;
      6: stateTransition = 11'd233;
      7: stateTransition = 11'd233;
      8: stateTransition = 11'd233;
      9: stateTransition = 11'd233;
      10: stateTransition = 11'd233;
      11: stateTransition = 11'd233;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd233;
      14: stateTransition = 11'd233;
      15: stateTransition = 11'd233;
      16: stateTransition = 11'd233;
      default: stateTransition = 11'bX;
    endcase
    234: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd234;
      2: stateTransition = 11'd234;
      3: stateTransition = 11'd234;
      4: stateTransition = 11'd234;
      5: stateTransition = 11'd234;
      6: stateTransition = 11'd234;
      7: stateTransition = 11'd234;
      8: stateTransition = 11'd234;
      9: stateTransition = 11'd234;
      10: stateTransition = 11'd234;
      11: stateTransition = 11'd234;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd234;
      14: stateTransition = 11'd234;
      15: stateTransition = 11'd234;
      16: stateTransition = 11'd234;
      default: stateTransition = 11'bX;
    endcase
    235: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd235;
      2: stateTransition = 11'd235;
      3: stateTransition = 11'd235;
      4: stateTransition = 11'd235;
      5: stateTransition = 11'd235;
      6: stateTransition = 11'd235;
      7: stateTransition = 11'd235;
      8: stateTransition = 11'd235;
      9: stateTransition = 11'd235;
      10: stateTransition = 11'd235;
      11: stateTransition = 11'd235;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd235;
      14: stateTransition = 11'd235;
      15: stateTransition = 11'd235;
      16: stateTransition = 11'd235;
      default: stateTransition = 11'bX;
    endcase
    236: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd236;
      2: stateTransition = 11'd236;
      3: stateTransition = 11'd236;
      4: stateTransition = 11'd236;
      5: stateTransition = 11'd236;
      6: stateTransition = 11'd236;
      7: stateTransition = 11'd236;
      8: stateTransition = 11'd236;
      9: stateTransition = 11'd236;
      10: stateTransition = 11'd236;
      11: stateTransition = 11'd236;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd236;
      14: stateTransition = 11'd236;
      15: stateTransition = 11'd236;
      16: stateTransition = 11'd236;
      default: stateTransition = 11'bX;
    endcase
    237: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd237;
      2: stateTransition = 11'd237;
      3: stateTransition = 11'd237;
      4: stateTransition = 11'd237;
      5: stateTransition = 11'd237;
      6: stateTransition = 11'd237;
      7: stateTransition = 11'd237;
      8: stateTransition = 11'd237;
      9: stateTransition = 11'd237;
      10: stateTransition = 11'd237;
      11: stateTransition = 11'd237;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd237;
      14: stateTransition = 11'd237;
      15: stateTransition = 11'd237;
      16: stateTransition = 11'd237;
      default: stateTransition = 11'bX;
    endcase
    238: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    239: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd239;
      2: stateTransition = 11'd239;
      3: stateTransition = 11'd239;
      4: stateTransition = 11'd239;
      5: stateTransition = 11'd239;
      6: stateTransition = 11'd239;
      7: stateTransition = 11'd239;
      8: stateTransition = 11'd239;
      9: stateTransition = 11'd239;
      10: stateTransition = 11'd239;
      11: stateTransition = 11'd239;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd239;
      14: stateTransition = 11'd239;
      15: stateTransition = 11'd239;
      16: stateTransition = 11'd239;
      default: stateTransition = 11'bX;
    endcase
    240: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd240;
      2: stateTransition = 11'd240;
      3: stateTransition = 11'd240;
      4: stateTransition = 11'd240;
      5: stateTransition = 11'd240;
      6: stateTransition = 11'd240;
      7: stateTransition = 11'd240;
      8: stateTransition = 11'd240;
      9: stateTransition = 11'd240;
      10: stateTransition = 11'd240;
      11: stateTransition = 11'd240;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd240;
      14: stateTransition = 11'd240;
      15: stateTransition = 11'd240;
      16: stateTransition = 11'd240;
      default: stateTransition = 11'bX;
    endcase
    241: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd241;
      2: stateTransition = 11'd241;
      3: stateTransition = 11'd241;
      4: stateTransition = 11'd241;
      5: stateTransition = 11'd241;
      6: stateTransition = 11'd241;
      7: stateTransition = 11'd241;
      8: stateTransition = 11'd241;
      9: stateTransition = 11'd241;
      10: stateTransition = 11'd241;
      11: stateTransition = 11'd241;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd241;
      14: stateTransition = 11'd241;
      15: stateTransition = 11'd241;
      16: stateTransition = 11'd241;
      default: stateTransition = 11'bX;
    endcase
    242: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd242;
      2: stateTransition = 11'd242;
      3: stateTransition = 11'd242;
      4: stateTransition = 11'd242;
      5: stateTransition = 11'd242;
      6: stateTransition = 11'd242;
      7: stateTransition = 11'd242;
      8: stateTransition = 11'd242;
      9: stateTransition = 11'd242;
      10: stateTransition = 11'd242;
      11: stateTransition = 11'd242;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd242;
      14: stateTransition = 11'd242;
      15: stateTransition = 11'd242;
      16: stateTransition = 11'd242;
      default: stateTransition = 11'bX;
    endcase
    243: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd243;
      2: stateTransition = 11'd243;
      3: stateTransition = 11'd243;
      4: stateTransition = 11'd243;
      5: stateTransition = 11'd243;
      6: stateTransition = 11'd243;
      7: stateTransition = 11'd243;
      8: stateTransition = 11'd243;
      9: stateTransition = 11'd243;
      10: stateTransition = 11'd243;
      11: stateTransition = 11'd243;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd243;
      14: stateTransition = 11'd243;
      15: stateTransition = 11'd243;
      16: stateTransition = 11'd243;
      default: stateTransition = 11'bX;
    endcase
    244: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd244;
      2: stateTransition = 11'd244;
      3: stateTransition = 11'd244;
      4: stateTransition = 11'd244;
      5: stateTransition = 11'd244;
      6: stateTransition = 11'd244;
      7: stateTransition = 11'd244;
      8: stateTransition = 11'd244;
      9: stateTransition = 11'd244;
      10: stateTransition = 11'd244;
      11: stateTransition = 11'd244;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd244;
      14: stateTransition = 11'd244;
      15: stateTransition = 11'd244;
      16: stateTransition = 11'd244;
      default: stateTransition = 11'bX;
    endcase
    245: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd245;
      2: stateTransition = 11'd245;
      3: stateTransition = 11'd245;
      4: stateTransition = 11'd245;
      5: stateTransition = 11'd245;
      6: stateTransition = 11'd245;
      7: stateTransition = 11'd245;
      8: stateTransition = 11'd245;
      9: stateTransition = 11'd245;
      10: stateTransition = 11'd245;
      11: stateTransition = 11'd245;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd245;
      14: stateTransition = 11'd245;
      15: stateTransition = 11'd245;
      16: stateTransition = 11'd245;
      default: stateTransition = 11'bX;
    endcase
    246: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd246;
      2: stateTransition = 11'd246;
      3: stateTransition = 11'd246;
      4: stateTransition = 11'd246;
      5: stateTransition = 11'd246;
      6: stateTransition = 11'd246;
      7: stateTransition = 11'd246;
      8: stateTransition = 11'd246;
      9: stateTransition = 11'd246;
      10: stateTransition = 11'd246;
      11: stateTransition = 11'd246;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd246;
      14: stateTransition = 11'd246;
      15: stateTransition = 11'd246;
      16: stateTransition = 11'd246;
      default: stateTransition = 11'bX;
    endcase
    247: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd247;
      2: stateTransition = 11'd247;
      3: stateTransition = 11'd247;
      4: stateTransition = 11'd247;
      5: stateTransition = 11'd247;
      6: stateTransition = 11'd247;
      7: stateTransition = 11'd247;
      8: stateTransition = 11'd247;
      9: stateTransition = 11'd247;
      10: stateTransition = 11'd247;
      11: stateTransition = 11'd247;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd247;
      14: stateTransition = 11'd247;
      15: stateTransition = 11'd247;
      16: stateTransition = 11'd247;
      default: stateTransition = 11'bX;
    endcase
    248: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd248;
      2: stateTransition = 11'd248;
      3: stateTransition = 11'd248;
      4: stateTransition = 11'd248;
      5: stateTransition = 11'd248;
      6: stateTransition = 11'd248;
      7: stateTransition = 11'd248;
      8: stateTransition = 11'd248;
      9: stateTransition = 11'd248;
      10: stateTransition = 11'd248;
      11: stateTransition = 11'd248;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd248;
      14: stateTransition = 11'd248;
      15: stateTransition = 11'd248;
      16: stateTransition = 11'd248;
      default: stateTransition = 11'bX;
    endcase
    249: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd249;
      2: stateTransition = 11'd249;
      3: stateTransition = 11'd249;
      4: stateTransition = 11'd249;
      5: stateTransition = 11'd249;
      6: stateTransition = 11'd249;
      7: stateTransition = 11'd249;
      8: stateTransition = 11'd249;
      9: stateTransition = 11'd249;
      10: stateTransition = 11'd249;
      11: stateTransition = 11'd249;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd249;
      14: stateTransition = 11'd249;
      15: stateTransition = 11'd249;
      16: stateTransition = 11'd249;
      default: stateTransition = 11'bX;
    endcase
    250: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd250;
      2: stateTransition = 11'd250;
      3: stateTransition = 11'd250;
      4: stateTransition = 11'd250;
      5: stateTransition = 11'd250;
      6: stateTransition = 11'd250;
      7: stateTransition = 11'd250;
      8: stateTransition = 11'd250;
      9: stateTransition = 11'd250;
      10: stateTransition = 11'd250;
      11: stateTransition = 11'd250;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd250;
      14: stateTransition = 11'd250;
      15: stateTransition = 11'd250;
      16: stateTransition = 11'd250;
      default: stateTransition = 11'bX;
    endcase
    251: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd251;
      2: stateTransition = 11'd251;
      3: stateTransition = 11'd251;
      4: stateTransition = 11'd251;
      5: stateTransition = 11'd251;
      6: stateTransition = 11'd251;
      7: stateTransition = 11'd251;
      8: stateTransition = 11'd251;
      9: stateTransition = 11'd251;
      10: stateTransition = 11'd251;
      11: stateTransition = 11'd251;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd251;
      14: stateTransition = 11'd251;
      15: stateTransition = 11'd251;
      16: stateTransition = 11'd251;
      default: stateTransition = 11'bX;
    endcase
    252: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd252;
      2: stateTransition = 11'd252;
      3: stateTransition = 11'd252;
      4: stateTransition = 11'd252;
      5: stateTransition = 11'd252;
      6: stateTransition = 11'd252;
      7: stateTransition = 11'd252;
      8: stateTransition = 11'd252;
      9: stateTransition = 11'd252;
      10: stateTransition = 11'd252;
      11: stateTransition = 11'd252;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd252;
      14: stateTransition = 11'd252;
      15: stateTransition = 11'd252;
      16: stateTransition = 11'd252;
      default: stateTransition = 11'bX;
    endcase
    253: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd253;
      2: stateTransition = 11'd253;
      3: stateTransition = 11'd253;
      4: stateTransition = 11'd253;
      5: stateTransition = 11'd253;
      6: stateTransition = 11'd253;
      7: stateTransition = 11'd253;
      8: stateTransition = 11'd253;
      9: stateTransition = 11'd253;
      10: stateTransition = 11'd253;
      11: stateTransition = 11'd253;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd253;
      14: stateTransition = 11'd253;
      15: stateTransition = 11'd253;
      16: stateTransition = 11'd253;
      default: stateTransition = 11'bX;
    endcase
    254: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd254;
      2: stateTransition = 11'd254;
      3: stateTransition = 11'd254;
      4: stateTransition = 11'd254;
      5: stateTransition = 11'd254;
      6: stateTransition = 11'd254;
      7: stateTransition = 11'd254;
      8: stateTransition = 11'd254;
      9: stateTransition = 11'd254;
      10: stateTransition = 11'd254;
      11: stateTransition = 11'd254;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd254;
      14: stateTransition = 11'd254;
      15: stateTransition = 11'd254;
      16: stateTransition = 11'd254;
      default: stateTransition = 11'bX;
    endcase
    255: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd255;
      2: stateTransition = 11'd255;
      3: stateTransition = 11'd255;
      4: stateTransition = 11'd255;
      5: stateTransition = 11'd255;
      6: stateTransition = 11'd255;
      7: stateTransition = 11'd255;
      8: stateTransition = 11'd255;
      9: stateTransition = 11'd255;
      10: stateTransition = 11'd255;
      11: stateTransition = 11'd255;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd255;
      14: stateTransition = 11'd255;
      15: stateTransition = 11'd255;
      16: stateTransition = 11'd255;
      default: stateTransition = 11'bX;
    endcase
    256: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd256;
      2: stateTransition = 11'd256;
      3: stateTransition = 11'd256;
      4: stateTransition = 11'd256;
      5: stateTransition = 11'd256;
      6: stateTransition = 11'd256;
      7: stateTransition = 11'd256;
      8: stateTransition = 11'd256;
      9: stateTransition = 11'd256;
      10: stateTransition = 11'd256;
      11: stateTransition = 11'd256;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd256;
      14: stateTransition = 11'd256;
      15: stateTransition = 11'd256;
      16: stateTransition = 11'd256;
      default: stateTransition = 11'bX;
    endcase
    257: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd257;
      2: stateTransition = 11'd257;
      3: stateTransition = 11'd257;
      4: stateTransition = 11'd257;
      5: stateTransition = 11'd257;
      6: stateTransition = 11'd257;
      7: stateTransition = 11'd257;
      8: stateTransition = 11'd257;
      9: stateTransition = 11'd257;
      10: stateTransition = 11'd257;
      11: stateTransition = 11'd257;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd257;
      14: stateTransition = 11'd257;
      15: stateTransition = 11'd257;
      16: stateTransition = 11'd257;
      default: stateTransition = 11'bX;
    endcase
    258: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd258;
      2: stateTransition = 11'd258;
      3: stateTransition = 11'd258;
      4: stateTransition = 11'd258;
      5: stateTransition = 11'd258;
      6: stateTransition = 11'd258;
      7: stateTransition = 11'd258;
      8: stateTransition = 11'd258;
      9: stateTransition = 11'd258;
      10: stateTransition = 11'd258;
      11: stateTransition = 11'd258;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd258;
      14: stateTransition = 11'd258;
      15: stateTransition = 11'd258;
      16: stateTransition = 11'd258;
      default: stateTransition = 11'bX;
    endcase
    259: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd259;
      2: stateTransition = 11'd259;
      3: stateTransition = 11'd259;
      4: stateTransition = 11'd259;
      5: stateTransition = 11'd259;
      6: stateTransition = 11'd259;
      7: stateTransition = 11'd259;
      8: stateTransition = 11'd259;
      9: stateTransition = 11'd259;
      10: stateTransition = 11'd259;
      11: stateTransition = 11'd259;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd259;
      14: stateTransition = 11'd259;
      15: stateTransition = 11'd259;
      16: stateTransition = 11'd259;
      default: stateTransition = 11'bX;
    endcase
    260: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd260;
      2: stateTransition = 11'd260;
      3: stateTransition = 11'd260;
      4: stateTransition = 11'd260;
      5: stateTransition = 11'd260;
      6: stateTransition = 11'd260;
      7: stateTransition = 11'd260;
      8: stateTransition = 11'd260;
      9: stateTransition = 11'd260;
      10: stateTransition = 11'd260;
      11: stateTransition = 11'd260;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd260;
      14: stateTransition = 11'd260;
      15: stateTransition = 11'd260;
      16: stateTransition = 11'd260;
      default: stateTransition = 11'bX;
    endcase
    261: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd261;
      2: stateTransition = 11'd261;
      3: stateTransition = 11'd261;
      4: stateTransition = 11'd261;
      5: stateTransition = 11'd261;
      6: stateTransition = 11'd261;
      7: stateTransition = 11'd261;
      8: stateTransition = 11'd261;
      9: stateTransition = 11'd261;
      10: stateTransition = 11'd261;
      11: stateTransition = 11'd261;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd261;
      14: stateTransition = 11'd261;
      15: stateTransition = 11'd261;
      16: stateTransition = 11'd261;
      default: stateTransition = 11'bX;
    endcase
    262: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd262;
      2: stateTransition = 11'd262;
      3: stateTransition = 11'd262;
      4: stateTransition = 11'd262;
      5: stateTransition = 11'd262;
      6: stateTransition = 11'd262;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd262;
      10: stateTransition = 11'd262;
      11: stateTransition = 11'd262;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd262;
      14: stateTransition = 11'd262;
      15: stateTransition = 11'd262;
      16: stateTransition = 11'd262;
      default: stateTransition = 11'bX;
    endcase
    263: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd263;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd263;
      4: stateTransition = 11'd263;
      5: stateTransition = 11'd263;
      6: stateTransition = 11'd263;
      7: stateTransition = 11'd263;
      8: stateTransition = 11'd263;
      9: stateTransition = 11'd263;
      10: stateTransition = 11'd263;
      11: stateTransition = 11'd263;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd263;
      14: stateTransition = 11'd263;
      15: stateTransition = 11'd263;
      16: stateTransition = 11'd263;
      default: stateTransition = 11'bX;
    endcase
    264: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd264;
      2: stateTransition = 11'd264;
      3: stateTransition = 11'd264;
      4: stateTransition = 11'd264;
      5: stateTransition = 11'd264;
      6: stateTransition = 11'd264;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd264;
      10: stateTransition = 11'd264;
      11: stateTransition = 11'd264;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd264;
      14: stateTransition = 11'd264;
      15: stateTransition = 11'd264;
      16: stateTransition = 11'd264;
      default: stateTransition = 11'bX;
    endcase
    265: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd265;
      2: stateTransition = 11'd265;
      3: stateTransition = 11'd265;
      4: stateTransition = 11'd265;
      5: stateTransition = 11'd265;
      6: stateTransition = 11'd265;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd265;
      10: stateTransition = 11'd265;
      11: stateTransition = 11'd265;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd265;
      14: stateTransition = 11'd265;
      15: stateTransition = 11'd265;
      16: stateTransition = 11'd265;
      default: stateTransition = 11'bX;
    endcase
    266: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd266;
      2: stateTransition = 11'd266;
      3: stateTransition = 11'd266;
      4: stateTransition = 11'd266;
      5: stateTransition = 11'd266;
      6: stateTransition = 11'd266;
      7: stateTransition = 11'd266;
      8: stateTransition = 11'd266;
      9: stateTransition = 11'd266;
      10: stateTransition = 11'd266;
      11: stateTransition = 11'd266;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd266;
      14: stateTransition = 11'd266;
      15: stateTransition = 11'd266;
      16: stateTransition = 11'd266;
      default: stateTransition = 11'bX;
    endcase
    267: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd267;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd267;
      4: stateTransition = 11'd267;
      5: stateTransition = 11'd267;
      6: stateTransition = 11'd267;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd267;
      9: stateTransition = 11'd267;
      10: stateTransition = 11'd267;
      11: stateTransition = 11'd267;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd267;
      14: stateTransition = 11'd267;
      15: stateTransition = 11'd267;
      16: stateTransition = 11'd267;
      default: stateTransition = 11'bX;
    endcase
    268: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd268;
      2: stateTransition = 11'd268;
      3: stateTransition = 11'd268;
      4: stateTransition = 11'd268;
      5: stateTransition = 11'd268;
      6: stateTransition = 11'd268;
      7: stateTransition = 11'd268;
      8: stateTransition = 11'd268;
      9: stateTransition = 11'd268;
      10: stateTransition = 11'd268;
      11: stateTransition = 11'd268;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd268;
      14: stateTransition = 11'd268;
      15: stateTransition = 11'd268;
      16: stateTransition = 11'd268;
      default: stateTransition = 11'bX;
    endcase
    269: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd269;
      2: stateTransition = 11'd269;
      3: stateTransition = 11'd269;
      4: stateTransition = 11'd269;
      5: stateTransition = 11'd269;
      6: stateTransition = 11'd269;
      7: stateTransition = 11'd269;
      8: stateTransition = 11'd269;
      9: stateTransition = 11'd269;
      10: stateTransition = 11'd269;
      11: stateTransition = 11'd269;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd269;
      14: stateTransition = 11'd269;
      15: stateTransition = 11'd269;
      16: stateTransition = 11'd269;
      default: stateTransition = 11'bX;
    endcase
    270: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd270;
      2: stateTransition = 11'd270;
      3: stateTransition = 11'd270;
      4: stateTransition = 11'd270;
      5: stateTransition = 11'd270;
      6: stateTransition = 11'd270;
      7: stateTransition = 11'd270;
      8: stateTransition = 11'd270;
      9: stateTransition = 11'd270;
      10: stateTransition = 11'd270;
      11: stateTransition = 11'd270;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd270;
      14: stateTransition = 11'd270;
      15: stateTransition = 11'd270;
      16: stateTransition = 11'd270;
      default: stateTransition = 11'bX;
    endcase
    271: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd271;
      2: stateTransition = 11'd271;
      3: stateTransition = 11'd271;
      4: stateTransition = 11'd271;
      5: stateTransition = 11'd271;
      6: stateTransition = 11'd271;
      7: stateTransition = 11'd271;
      8: stateTransition = 11'd271;
      9: stateTransition = 11'd271;
      10: stateTransition = 11'd271;
      11: stateTransition = 11'd271;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd271;
      14: stateTransition = 11'd271;
      15: stateTransition = 11'd271;
      16: stateTransition = 11'd271;
      default: stateTransition = 11'bX;
    endcase
    272: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd272;
      2: stateTransition = 11'd272;
      3: stateTransition = 11'd272;
      4: stateTransition = 11'd272;
      5: stateTransition = 11'd272;
      6: stateTransition = 11'd272;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd272;
      10: stateTransition = 11'd272;
      11: stateTransition = 11'd272;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd272;
      14: stateTransition = 11'd272;
      15: stateTransition = 11'd272;
      16: stateTransition = 11'd272;
      default: stateTransition = 11'bX;
    endcase
    273: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd273;
      2: stateTransition = 11'd273;
      3: stateTransition = 11'd273;
      4: stateTransition = 11'd273;
      5: stateTransition = 11'd273;
      6: stateTransition = 11'd273;
      7: stateTransition = 11'd273;
      8: stateTransition = 11'd273;
      9: stateTransition = 11'd273;
      10: stateTransition = 11'd273;
      11: stateTransition = 11'd273;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd273;
      14: stateTransition = 11'd273;
      15: stateTransition = 11'd273;
      16: stateTransition = 11'd273;
      default: stateTransition = 11'bX;
    endcase
    274: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    275: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd275;
      2: stateTransition = 11'd275;
      3: stateTransition = 11'd275;
      4: stateTransition = 11'd275;
      5: stateTransition = 11'd275;
      6: stateTransition = 11'd275;
      7: stateTransition = 11'd275;
      8: stateTransition = 11'd275;
      9: stateTransition = 11'd275;
      10: stateTransition = 11'd275;
      11: stateTransition = 11'd275;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd275;
      14: stateTransition = 11'd275;
      15: stateTransition = 11'd275;
      16: stateTransition = 11'd275;
      default: stateTransition = 11'bX;
    endcase
    276: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd276;
      2: stateTransition = 11'd276;
      3: stateTransition = 11'd276;
      4: stateTransition = 11'd276;
      5: stateTransition = 11'd276;
      6: stateTransition = 11'd276;
      7: stateTransition = 11'd276;
      8: stateTransition = 11'd276;
      9: stateTransition = 11'd276;
      10: stateTransition = 11'd276;
      11: stateTransition = 11'd276;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd276;
      14: stateTransition = 11'd276;
      15: stateTransition = 11'd276;
      16: stateTransition = 11'd276;
      default: stateTransition = 11'bX;
    endcase
    277: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd277;
      2: stateTransition = 11'd277;
      3: stateTransition = 11'd277;
      4: stateTransition = 11'd277;
      5: stateTransition = 11'd277;
      6: stateTransition = 11'd277;
      7: stateTransition = 11'd277;
      8: stateTransition = 11'd277;
      9: stateTransition = 11'd277;
      10: stateTransition = 11'd277;
      11: stateTransition = 11'd277;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd277;
      14: stateTransition = 11'd277;
      15: stateTransition = 11'd277;
      16: stateTransition = 11'd277;
      default: stateTransition = 11'bX;
    endcase
    278: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd278;
      2: stateTransition = 11'd278;
      3: stateTransition = 11'd278;
      4: stateTransition = 11'd278;
      5: stateTransition = 11'd278;
      6: stateTransition = 11'd278;
      7: stateTransition = 11'd278;
      8: stateTransition = 11'd278;
      9: stateTransition = 11'd278;
      10: stateTransition = 11'd278;
      11: stateTransition = 11'd278;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd278;
      14: stateTransition = 11'd278;
      15: stateTransition = 11'd278;
      16: stateTransition = 11'd278;
      default: stateTransition = 11'bX;
    endcase
    279: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd279;
      2: stateTransition = 11'd279;
      3: stateTransition = 11'd279;
      4: stateTransition = 11'd279;
      5: stateTransition = 11'd279;
      6: stateTransition = 11'd279;
      7: stateTransition = 11'd279;
      8: stateTransition = 11'd279;
      9: stateTransition = 11'd279;
      10: stateTransition = 11'd279;
      11: stateTransition = 11'd279;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd279;
      14: stateTransition = 11'd279;
      15: stateTransition = 11'd279;
      16: stateTransition = 11'd279;
      default: stateTransition = 11'bX;
    endcase
    280: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd280;
      2: stateTransition = 11'd280;
      3: stateTransition = 11'd280;
      4: stateTransition = 11'd280;
      5: stateTransition = 11'd280;
      6: stateTransition = 11'd280;
      7: stateTransition = 11'd280;
      8: stateTransition = 11'd280;
      9: stateTransition = 11'd280;
      10: stateTransition = 11'd280;
      11: stateTransition = 11'd280;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd280;
      14: stateTransition = 11'd280;
      15: stateTransition = 11'd280;
      16: stateTransition = 11'd280;
      default: stateTransition = 11'bX;
    endcase
    281: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd281;
      2: stateTransition = 11'd281;
      3: stateTransition = 11'd281;
      4: stateTransition = 11'd281;
      5: stateTransition = 11'd281;
      6: stateTransition = 11'd281;
      7: stateTransition = 11'd281;
      8: stateTransition = 11'd281;
      9: stateTransition = 11'd281;
      10: stateTransition = 11'd281;
      11: stateTransition = 11'd281;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd281;
      14: stateTransition = 11'd281;
      15: stateTransition = 11'd281;
      16: stateTransition = 11'd281;
      default: stateTransition = 11'bX;
    endcase
    282: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd282;
      2: stateTransition = 11'd282;
      3: stateTransition = 11'd282;
      4: stateTransition = 11'd282;
      5: stateTransition = 11'd282;
      6: stateTransition = 11'd282;
      7: stateTransition = 11'd282;
      8: stateTransition = 11'd282;
      9: stateTransition = 11'd282;
      10: stateTransition = 11'd282;
      11: stateTransition = 11'd282;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd282;
      14: stateTransition = 11'd282;
      15: stateTransition = 11'd282;
      16: stateTransition = 11'd282;
      default: stateTransition = 11'bX;
    endcase
    283: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd283;
      2: stateTransition = 11'd283;
      3: stateTransition = 11'd283;
      4: stateTransition = 11'd283;
      5: stateTransition = 11'd283;
      6: stateTransition = 11'd283;
      7: stateTransition = 11'd283;
      8: stateTransition = 11'd283;
      9: stateTransition = 11'd283;
      10: stateTransition = 11'd283;
      11: stateTransition = 11'd283;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd283;
      14: stateTransition = 11'd283;
      15: stateTransition = 11'd283;
      16: stateTransition = 11'd283;
      default: stateTransition = 11'bX;
    endcase
    284: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd284;
      2: stateTransition = 11'd284;
      3: stateTransition = 11'd284;
      4: stateTransition = 11'd284;
      5: stateTransition = 11'd284;
      6: stateTransition = 11'd284;
      7: stateTransition = 11'd284;
      8: stateTransition = 11'd284;
      9: stateTransition = 11'd284;
      10: stateTransition = 11'd284;
      11: stateTransition = 11'd284;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd284;
      14: stateTransition = 11'd284;
      15: stateTransition = 11'd284;
      16: stateTransition = 11'd284;
      default: stateTransition = 11'bX;
    endcase
    285: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd285;
      2: stateTransition = 11'd285;
      3: stateTransition = 11'd285;
      4: stateTransition = 11'd285;
      5: stateTransition = 11'd285;
      6: stateTransition = 11'd285;
      7: stateTransition = 11'd285;
      8: stateTransition = 11'd285;
      9: stateTransition = 11'd285;
      10: stateTransition = 11'd285;
      11: stateTransition = 11'd285;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd285;
      14: stateTransition = 11'd285;
      15: stateTransition = 11'd285;
      16: stateTransition = 11'd285;
      default: stateTransition = 11'bX;
    endcase
    286: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd286;
      2: stateTransition = 11'd286;
      3: stateTransition = 11'd286;
      4: stateTransition = 11'd286;
      5: stateTransition = 11'd286;
      6: stateTransition = 11'd286;
      7: stateTransition = 11'd286;
      8: stateTransition = 11'd286;
      9: stateTransition = 11'd286;
      10: stateTransition = 11'd286;
      11: stateTransition = 11'd286;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd286;
      14: stateTransition = 11'd286;
      15: stateTransition = 11'd286;
      16: stateTransition = 11'd286;
      default: stateTransition = 11'bX;
    endcase
    287: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd287;
      2: stateTransition = 11'd287;
      3: stateTransition = 11'd287;
      4: stateTransition = 11'd287;
      5: stateTransition = 11'd287;
      6: stateTransition = 11'd287;
      7: stateTransition = 11'd287;
      8: stateTransition = 11'd287;
      9: stateTransition = 11'd287;
      10: stateTransition = 11'd287;
      11: stateTransition = 11'd287;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd287;
      14: stateTransition = 11'd287;
      15: stateTransition = 11'd287;
      16: stateTransition = 11'd287;
      default: stateTransition = 11'bX;
    endcase
    288: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd288;
      2: stateTransition = 11'd288;
      3: stateTransition = 11'd288;
      4: stateTransition = 11'd288;
      5: stateTransition = 11'd288;
      6: stateTransition = 11'd288;
      7: stateTransition = 11'd288;
      8: stateTransition = 11'd288;
      9: stateTransition = 11'd288;
      10: stateTransition = 11'd288;
      11: stateTransition = 11'd288;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd288;
      14: stateTransition = 11'd288;
      15: stateTransition = 11'd288;
      16: stateTransition = 11'd288;
      default: stateTransition = 11'bX;
    endcase
    289: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd289;
      2: stateTransition = 11'd289;
      3: stateTransition = 11'd289;
      4: stateTransition = 11'd289;
      5: stateTransition = 11'd289;
      6: stateTransition = 11'd289;
      7: stateTransition = 11'd289;
      8: stateTransition = 11'd289;
      9: stateTransition = 11'd289;
      10: stateTransition = 11'd289;
      11: stateTransition = 11'd289;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd289;
      14: stateTransition = 11'd289;
      15: stateTransition = 11'd289;
      16: stateTransition = 11'd289;
      default: stateTransition = 11'bX;
    endcase
    290: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd290;
      2: stateTransition = 11'd290;
      3: stateTransition = 11'd290;
      4: stateTransition = 11'd290;
      5: stateTransition = 11'd290;
      6: stateTransition = 11'd290;
      7: stateTransition = 11'd290;
      8: stateTransition = 11'd290;
      9: stateTransition = 11'd290;
      10: stateTransition = 11'd290;
      11: stateTransition = 11'd290;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd290;
      14: stateTransition = 11'd290;
      15: stateTransition = 11'd290;
      16: stateTransition = 11'd290;
      default: stateTransition = 11'bX;
    endcase
    291: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd291;
      2: stateTransition = 11'd291;
      3: stateTransition = 11'd291;
      4: stateTransition = 11'd291;
      5: stateTransition = 11'd291;
      6: stateTransition = 11'd291;
      7: stateTransition = 11'd291;
      8: stateTransition = 11'd291;
      9: stateTransition = 11'd291;
      10: stateTransition = 11'd291;
      11: stateTransition = 11'd291;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd291;
      14: stateTransition = 11'd291;
      15: stateTransition = 11'd291;
      16: stateTransition = 11'd291;
      default: stateTransition = 11'bX;
    endcase
    292: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd292;
      2: stateTransition = 11'd292;
      3: stateTransition = 11'd292;
      4: stateTransition = 11'd292;
      5: stateTransition = 11'd292;
      6: stateTransition = 11'd292;
      7: stateTransition = 11'd292;
      8: stateTransition = 11'd292;
      9: stateTransition = 11'd292;
      10: stateTransition = 11'd292;
      11: stateTransition = 11'd292;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd292;
      14: stateTransition = 11'd292;
      15: stateTransition = 11'd292;
      16: stateTransition = 11'd292;
      default: stateTransition = 11'bX;
    endcase
    293: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd293;
      2: stateTransition = 11'd293;
      3: stateTransition = 11'd293;
      4: stateTransition = 11'd293;
      5: stateTransition = 11'd293;
      6: stateTransition = 11'd293;
      7: stateTransition = 11'd293;
      8: stateTransition = 11'd293;
      9: stateTransition = 11'd293;
      10: stateTransition = 11'd293;
      11: stateTransition = 11'd293;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd293;
      14: stateTransition = 11'd293;
      15: stateTransition = 11'd293;
      16: stateTransition = 11'd293;
      default: stateTransition = 11'bX;
    endcase
    294: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd294;
      2: stateTransition = 11'd294;
      3: stateTransition = 11'd294;
      4: stateTransition = 11'd294;
      5: stateTransition = 11'd294;
      6: stateTransition = 11'd294;
      7: stateTransition = 11'd294;
      8: stateTransition = 11'd294;
      9: stateTransition = 11'd294;
      10: stateTransition = 11'd294;
      11: stateTransition = 11'd294;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd294;
      14: stateTransition = 11'd294;
      15: stateTransition = 11'd294;
      16: stateTransition = 11'd294;
      default: stateTransition = 11'bX;
    endcase
    295: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd295;
      2: stateTransition = 11'd295;
      3: stateTransition = 11'd295;
      4: stateTransition = 11'd295;
      5: stateTransition = 11'd295;
      6: stateTransition = 11'd295;
      7: stateTransition = 11'd295;
      8: stateTransition = 11'd295;
      9: stateTransition = 11'd295;
      10: stateTransition = 11'd295;
      11: stateTransition = 11'd295;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd295;
      14: stateTransition = 11'd295;
      15: stateTransition = 11'd295;
      16: stateTransition = 11'd295;
      default: stateTransition = 11'bX;
    endcase
    296: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd296;
      2: stateTransition = 11'd296;
      3: stateTransition = 11'd296;
      4: stateTransition = 11'd296;
      5: stateTransition = 11'd296;
      6: stateTransition = 11'd296;
      7: stateTransition = 11'd296;
      8: stateTransition = 11'd296;
      9: stateTransition = 11'd296;
      10: stateTransition = 11'd296;
      11: stateTransition = 11'd296;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd296;
      14: stateTransition = 11'd296;
      15: stateTransition = 11'd296;
      16: stateTransition = 11'd296;
      default: stateTransition = 11'bX;
    endcase
    297: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd297;
      2: stateTransition = 11'd297;
      3: stateTransition = 11'd297;
      4: stateTransition = 11'd297;
      5: stateTransition = 11'd297;
      6: stateTransition = 11'd297;
      7: stateTransition = 11'd297;
      8: stateTransition = 11'd297;
      9: stateTransition = 11'd297;
      10: stateTransition = 11'd297;
      11: stateTransition = 11'd297;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd297;
      14: stateTransition = 11'd297;
      15: stateTransition = 11'd297;
      16: stateTransition = 11'd297;
      default: stateTransition = 11'bX;
    endcase
    298: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd298;
      2: stateTransition = 11'd298;
      3: stateTransition = 11'd298;
      4: stateTransition = 11'd298;
      5: stateTransition = 11'd298;
      6: stateTransition = 11'd298;
      7: stateTransition = 11'd298;
      8: stateTransition = 11'd298;
      9: stateTransition = 11'd298;
      10: stateTransition = 11'd298;
      11: stateTransition = 11'd298;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd298;
      14: stateTransition = 11'd298;
      15: stateTransition = 11'd298;
      16: stateTransition = 11'd298;
      default: stateTransition = 11'bX;
    endcase
    299: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd299;
      2: stateTransition = 11'd299;
      3: stateTransition = 11'd299;
      4: stateTransition = 11'd299;
      5: stateTransition = 11'd299;
      6: stateTransition = 11'd299;
      7: stateTransition = 11'd299;
      8: stateTransition = 11'd299;
      9: stateTransition = 11'd299;
      10: stateTransition = 11'd299;
      11: stateTransition = 11'd299;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd299;
      14: stateTransition = 11'd299;
      15: stateTransition = 11'd299;
      16: stateTransition = 11'd299;
      default: stateTransition = 11'bX;
    endcase
    300: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd300;
      2: stateTransition = 11'd300;
      3: stateTransition = 11'd300;
      4: stateTransition = 11'd300;
      5: stateTransition = 11'd300;
      6: stateTransition = 11'd300;
      7: stateTransition = 11'd300;
      8: stateTransition = 11'd300;
      9: stateTransition = 11'd300;
      10: stateTransition = 11'd300;
      11: stateTransition = 11'd300;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd300;
      14: stateTransition = 11'd300;
      15: stateTransition = 11'd300;
      16: stateTransition = 11'd300;
      default: stateTransition = 11'bX;
    endcase
    301: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd301;
      2: stateTransition = 11'd301;
      3: stateTransition = 11'd301;
      4: stateTransition = 11'd301;
      5: stateTransition = 11'd301;
      6: stateTransition = 11'd301;
      7: stateTransition = 11'd301;
      8: stateTransition = 11'd301;
      9: stateTransition = 11'd301;
      10: stateTransition = 11'd301;
      11: stateTransition = 11'd301;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd301;
      14: stateTransition = 11'd301;
      15: stateTransition = 11'd301;
      16: stateTransition = 11'd301;
      default: stateTransition = 11'bX;
    endcase
    302: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd302;
      2: stateTransition = 11'd302;
      3: stateTransition = 11'd302;
      4: stateTransition = 11'd302;
      5: stateTransition = 11'd302;
      6: stateTransition = 11'd302;
      7: stateTransition = 11'd302;
      8: stateTransition = 11'd302;
      9: stateTransition = 11'd302;
      10: stateTransition = 11'd302;
      11: stateTransition = 11'd302;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd302;
      14: stateTransition = 11'd302;
      15: stateTransition = 11'd302;
      16: stateTransition = 11'd302;
      default: stateTransition = 11'bX;
    endcase
    303: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd303;
      2: stateTransition = 11'd303;
      3: stateTransition = 11'd303;
      4: stateTransition = 11'd303;
      5: stateTransition = 11'd303;
      6: stateTransition = 11'd303;
      7: stateTransition = 11'd303;
      8: stateTransition = 11'd303;
      9: stateTransition = 11'd303;
      10: stateTransition = 11'd303;
      11: stateTransition = 11'd303;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd303;
      14: stateTransition = 11'd303;
      15: stateTransition = 11'd303;
      16: stateTransition = 11'd303;
      default: stateTransition = 11'bX;
    endcase
    304: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd304;
      2: stateTransition = 11'd304;
      3: stateTransition = 11'd304;
      4: stateTransition = 11'd304;
      5: stateTransition = 11'd304;
      6: stateTransition = 11'd304;
      7: stateTransition = 11'd304;
      8: stateTransition = 11'd304;
      9: stateTransition = 11'd304;
      10: stateTransition = 11'd304;
      11: stateTransition = 11'd304;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd304;
      14: stateTransition = 11'd304;
      15: stateTransition = 11'd304;
      16: stateTransition = 11'd304;
      default: stateTransition = 11'bX;
    endcase
    305: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd305;
      2: stateTransition = 11'd305;
      3: stateTransition = 11'd305;
      4: stateTransition = 11'd305;
      5: stateTransition = 11'd305;
      6: stateTransition = 11'd305;
      7: stateTransition = 11'd305;
      8: stateTransition = 11'd305;
      9: stateTransition = 11'd305;
      10: stateTransition = 11'd305;
      11: stateTransition = 11'd305;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd305;
      14: stateTransition = 11'd305;
      15: stateTransition = 11'd305;
      16: stateTransition = 11'd305;
      default: stateTransition = 11'bX;
    endcase
    306: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd306;
      2: stateTransition = 11'd306;
      3: stateTransition = 11'd306;
      4: stateTransition = 11'd306;
      5: stateTransition = 11'd306;
      6: stateTransition = 11'd306;
      7: stateTransition = 11'd306;
      8: stateTransition = 11'd306;
      9: stateTransition = 11'd306;
      10: stateTransition = 11'd306;
      11: stateTransition = 11'd306;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd306;
      14: stateTransition = 11'd306;
      15: stateTransition = 11'd306;
      16: stateTransition = 11'd306;
      default: stateTransition = 11'bX;
    endcase
    307: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd307;
      2: stateTransition = 11'd307;
      3: stateTransition = 11'd307;
      4: stateTransition = 11'd307;
      5: stateTransition = 11'd307;
      6: stateTransition = 11'd307;
      7: stateTransition = 11'd307;
      8: stateTransition = 11'd307;
      9: stateTransition = 11'd307;
      10: stateTransition = 11'd307;
      11: stateTransition = 11'd307;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd307;
      14: stateTransition = 11'd307;
      15: stateTransition = 11'd307;
      16: stateTransition = 11'd307;
      default: stateTransition = 11'bX;
    endcase
    308: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd308;
      2: stateTransition = 11'd308;
      3: stateTransition = 11'd308;
      4: stateTransition = 11'd308;
      5: stateTransition = 11'd308;
      6: stateTransition = 11'd308;
      7: stateTransition = 11'd308;
      8: stateTransition = 11'd308;
      9: stateTransition = 11'd308;
      10: stateTransition = 11'd308;
      11: stateTransition = 11'd308;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd308;
      14: stateTransition = 11'd308;
      15: stateTransition = 11'd308;
      16: stateTransition = 11'd308;
      default: stateTransition = 11'bX;
    endcase
    309: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd309;
      2: stateTransition = 11'd309;
      3: stateTransition = 11'd309;
      4: stateTransition = 11'd309;
      5: stateTransition = 11'd309;
      6: stateTransition = 11'd309;
      7: stateTransition = 11'd309;
      8: stateTransition = 11'd309;
      9: stateTransition = 11'd309;
      10: stateTransition = 11'd309;
      11: stateTransition = 11'd309;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd309;
      14: stateTransition = 11'd309;
      15: stateTransition = 11'd309;
      16: stateTransition = 11'd309;
      default: stateTransition = 11'bX;
    endcase
    310: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd310;
      2: stateTransition = 11'd310;
      3: stateTransition = 11'd310;
      4: stateTransition = 11'd310;
      5: stateTransition = 11'd310;
      6: stateTransition = 11'd310;
      7: stateTransition = 11'd310;
      8: stateTransition = 11'd310;
      9: stateTransition = 11'd310;
      10: stateTransition = 11'd310;
      11: stateTransition = 11'd310;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd310;
      14: stateTransition = 11'd310;
      15: stateTransition = 11'd310;
      16: stateTransition = 11'd310;
      default: stateTransition = 11'bX;
    endcase
    311: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd311;
      2: stateTransition = 11'd311;
      3: stateTransition = 11'd311;
      4: stateTransition = 11'd311;
      5: stateTransition = 11'd311;
      6: stateTransition = 11'd311;
      7: stateTransition = 11'd311;
      8: stateTransition = 11'd311;
      9: stateTransition = 11'd311;
      10: stateTransition = 11'd311;
      11: stateTransition = 11'd311;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd311;
      14: stateTransition = 11'd311;
      15: stateTransition = 11'd311;
      16: stateTransition = 11'd311;
      default: stateTransition = 11'bX;
    endcase
    312: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd312;
      2: stateTransition = 11'd312;
      3: stateTransition = 11'd312;
      4: stateTransition = 11'd312;
      5: stateTransition = 11'd312;
      6: stateTransition = 11'd312;
      7: stateTransition = 11'd312;
      8: stateTransition = 11'd312;
      9: stateTransition = 11'd312;
      10: stateTransition = 11'd312;
      11: stateTransition = 11'd312;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd312;
      14: stateTransition = 11'd312;
      15: stateTransition = 11'd312;
      16: stateTransition = 11'd312;
      default: stateTransition = 11'bX;
    endcase
    313: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd313;
      2: stateTransition = 11'd313;
      3: stateTransition = 11'd313;
      4: stateTransition = 11'd313;
      5: stateTransition = 11'd313;
      6: stateTransition = 11'd313;
      7: stateTransition = 11'd313;
      8: stateTransition = 11'd313;
      9: stateTransition = 11'd313;
      10: stateTransition = 11'd313;
      11: stateTransition = 11'd313;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd313;
      14: stateTransition = 11'd313;
      15: stateTransition = 11'd313;
      16: stateTransition = 11'd313;
      default: stateTransition = 11'bX;
    endcase
    314: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd314;
      2: stateTransition = 11'd314;
      3: stateTransition = 11'd314;
      4: stateTransition = 11'd314;
      5: stateTransition = 11'd314;
      6: stateTransition = 11'd314;
      7: stateTransition = 11'd314;
      8: stateTransition = 11'd314;
      9: stateTransition = 11'd314;
      10: stateTransition = 11'd314;
      11: stateTransition = 11'd314;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd314;
      14: stateTransition = 11'd314;
      15: stateTransition = 11'd314;
      16: stateTransition = 11'd314;
      default: stateTransition = 11'bX;
    endcase
    315: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd315;
      2: stateTransition = 11'd315;
      3: stateTransition = 11'd315;
      4: stateTransition = 11'd315;
      5: stateTransition = 11'd315;
      6: stateTransition = 11'd315;
      7: stateTransition = 11'd315;
      8: stateTransition = 11'd315;
      9: stateTransition = 11'd315;
      10: stateTransition = 11'd315;
      11: stateTransition = 11'd315;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd315;
      14: stateTransition = 11'd315;
      15: stateTransition = 11'd315;
      16: stateTransition = 11'd315;
      default: stateTransition = 11'bX;
    endcase
    316: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    317: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd317;
      2: stateTransition = 11'd317;
      3: stateTransition = 11'd317;
      4: stateTransition = 11'd317;
      5: stateTransition = 11'd317;
      6: stateTransition = 11'd317;
      7: stateTransition = 11'd317;
      8: stateTransition = 11'd317;
      9: stateTransition = 11'd317;
      10: stateTransition = 11'd317;
      11: stateTransition = 11'd317;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd317;
      14: stateTransition = 11'd317;
      15: stateTransition = 11'd317;
      16: stateTransition = 11'd317;
      default: stateTransition = 11'bX;
    endcase
    318: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd318;
      2: stateTransition = 11'd318;
      3: stateTransition = 11'd318;
      4: stateTransition = 11'd318;
      5: stateTransition = 11'd318;
      6: stateTransition = 11'd318;
      7: stateTransition = 11'd318;
      8: stateTransition = 11'd318;
      9: stateTransition = 11'd318;
      10: stateTransition = 11'd318;
      11: stateTransition = 11'd318;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd318;
      14: stateTransition = 11'd318;
      15: stateTransition = 11'd318;
      16: stateTransition = 11'd318;
      default: stateTransition = 11'bX;
    endcase
    319: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd319;
      2: stateTransition = 11'd319;
      3: stateTransition = 11'd319;
      4: stateTransition = 11'd319;
      5: stateTransition = 11'd319;
      6: stateTransition = 11'd319;
      7: stateTransition = 11'd319;
      8: stateTransition = 11'd319;
      9: stateTransition = 11'd319;
      10: stateTransition = 11'd319;
      11: stateTransition = 11'd319;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd319;
      14: stateTransition = 11'd319;
      15: stateTransition = 11'd319;
      16: stateTransition = 11'd319;
      default: stateTransition = 11'bX;
    endcase
    320: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd320;
      2: stateTransition = 11'd320;
      3: stateTransition = 11'd320;
      4: stateTransition = 11'd320;
      5: stateTransition = 11'd320;
      6: stateTransition = 11'd320;
      7: stateTransition = 11'd320;
      8: stateTransition = 11'd320;
      9: stateTransition = 11'd320;
      10: stateTransition = 11'd320;
      11: stateTransition = 11'd320;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd320;
      14: stateTransition = 11'd320;
      15: stateTransition = 11'd320;
      16: stateTransition = 11'd320;
      default: stateTransition = 11'bX;
    endcase
    321: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd321;
      2: stateTransition = 11'd321;
      3: stateTransition = 11'd321;
      4: stateTransition = 11'd321;
      5: stateTransition = 11'd321;
      6: stateTransition = 11'd321;
      7: stateTransition = 11'd321;
      8: stateTransition = 11'd321;
      9: stateTransition = 11'd321;
      10: stateTransition = 11'd321;
      11: stateTransition = 11'd321;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd321;
      14: stateTransition = 11'd321;
      15: stateTransition = 11'd321;
      16: stateTransition = 11'd321;
      default: stateTransition = 11'bX;
    endcase
    322: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd322;
      2: stateTransition = 11'd322;
      3: stateTransition = 11'd322;
      4: stateTransition = 11'd322;
      5: stateTransition = 11'd322;
      6: stateTransition = 11'd322;
      7: stateTransition = 11'd322;
      8: stateTransition = 11'd322;
      9: stateTransition = 11'd322;
      10: stateTransition = 11'd322;
      11: stateTransition = 11'd322;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd322;
      14: stateTransition = 11'd322;
      15: stateTransition = 11'd322;
      16: stateTransition = 11'd322;
      default: stateTransition = 11'bX;
    endcase
    323: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd323;
      2: stateTransition = 11'd323;
      3: stateTransition = 11'd323;
      4: stateTransition = 11'd323;
      5: stateTransition = 11'd323;
      6: stateTransition = 11'd323;
      7: stateTransition = 11'd323;
      8: stateTransition = 11'd323;
      9: stateTransition = 11'd323;
      10: stateTransition = 11'd323;
      11: stateTransition = 11'd323;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd323;
      14: stateTransition = 11'd323;
      15: stateTransition = 11'd323;
      16: stateTransition = 11'd323;
      default: stateTransition = 11'bX;
    endcase
    324: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd324;
      2: stateTransition = 11'd324;
      3: stateTransition = 11'd324;
      4: stateTransition = 11'd324;
      5: stateTransition = 11'd324;
      6: stateTransition = 11'd324;
      7: stateTransition = 11'd324;
      8: stateTransition = 11'd324;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd324;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd324;
      default: stateTransition = 11'bX;
    endcase
    325: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd325;
      2: stateTransition = 11'd325;
      3: stateTransition = 11'd325;
      4: stateTransition = 11'd325;
      5: stateTransition = 11'd325;
      6: stateTransition = 11'd325;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd325;
      10: stateTransition = 11'd325;
      11: stateTransition = 11'd325;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd325;
      14: stateTransition = 11'd325;
      15: stateTransition = 11'd325;
      16: stateTransition = 11'd325;
      default: stateTransition = 11'bX;
    endcase
    326: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd326;
      2: stateTransition = 11'd326;
      3: stateTransition = 11'd326;
      4: stateTransition = 11'd326;
      5: stateTransition = 11'd326;
      6: stateTransition = 11'd326;
      7: stateTransition = 11'd326;
      8: stateTransition = 11'd326;
      9: stateTransition = 11'd326;
      10: stateTransition = 11'd326;
      11: stateTransition = 11'd326;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd326;
      14: stateTransition = 11'd326;
      15: stateTransition = 11'd326;
      16: stateTransition = 11'd326;
      default: stateTransition = 11'bX;
    endcase
    327: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd327;
      2: stateTransition = 11'd327;
      3: stateTransition = 11'd327;
      4: stateTransition = 11'd327;
      5: stateTransition = 11'd327;
      6: stateTransition = 11'd327;
      7: stateTransition = 11'd327;
      8: stateTransition = 11'd327;
      9: stateTransition = 11'd327;
      10: stateTransition = 11'd327;
      11: stateTransition = 11'd327;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd327;
      14: stateTransition = 11'd327;
      15: stateTransition = 11'd327;
      16: stateTransition = 11'd327;
      default: stateTransition = 11'bX;
    endcase
    328: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd328;
      2: stateTransition = 11'd328;
      3: stateTransition = 11'd328;
      4: stateTransition = 11'd328;
      5: stateTransition = 11'd328;
      6: stateTransition = 11'd328;
      7: stateTransition = 11'd328;
      8: stateTransition = 11'd328;
      9: stateTransition = 11'd328;
      10: stateTransition = 11'd328;
      11: stateTransition = 11'd328;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd328;
      14: stateTransition = 11'd328;
      15: stateTransition = 11'd328;
      16: stateTransition = 11'd328;
      default: stateTransition = 11'bX;
    endcase
    329: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd329;
      2: stateTransition = 11'd329;
      3: stateTransition = 11'd329;
      4: stateTransition = 11'd329;
      5: stateTransition = 11'd329;
      6: stateTransition = 11'd329;
      7: stateTransition = 11'd329;
      8: stateTransition = 11'd329;
      9: stateTransition = 11'd329;
      10: stateTransition = 11'd329;
      11: stateTransition = 11'd329;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd329;
      14: stateTransition = 11'd329;
      15: stateTransition = 11'd329;
      16: stateTransition = 11'd329;
      default: stateTransition = 11'bX;
    endcase
    330: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd330;
      2: stateTransition = 11'd330;
      3: stateTransition = 11'd330;
      4: stateTransition = 11'd330;
      5: stateTransition = 11'd330;
      6: stateTransition = 11'd330;
      7: stateTransition = 11'd330;
      8: stateTransition = 11'd330;
      9: stateTransition = 11'd330;
      10: stateTransition = 11'd330;
      11: stateTransition = 11'd330;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd330;
      14: stateTransition = 11'd330;
      15: stateTransition = 11'd330;
      16: stateTransition = 11'd330;
      default: stateTransition = 11'bX;
    endcase
    331: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd331;
      2: stateTransition = 11'd331;
      3: stateTransition = 11'd331;
      4: stateTransition = 11'd331;
      5: stateTransition = 11'd331;
      6: stateTransition = 11'd331;
      7: stateTransition = 11'd331;
      8: stateTransition = 11'd331;
      9: stateTransition = 11'd331;
      10: stateTransition = 11'd331;
      11: stateTransition = 11'd331;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd331;
      14: stateTransition = 11'd331;
      15: stateTransition = 11'd331;
      16: stateTransition = 11'd331;
      default: stateTransition = 11'bX;
    endcase
    332: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd332;
      2: stateTransition = 11'd332;
      3: stateTransition = 11'd332;
      4: stateTransition = 11'd332;
      5: stateTransition = 11'd332;
      6: stateTransition = 11'd332;
      7: stateTransition = 11'd332;
      8: stateTransition = 11'd332;
      9: stateTransition = 11'd332;
      10: stateTransition = 11'd332;
      11: stateTransition = 11'd332;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd332;
      14: stateTransition = 11'd332;
      15: stateTransition = 11'd332;
      16: stateTransition = 11'd332;
      default: stateTransition = 11'bX;
    endcase
    333: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd333;
      2: stateTransition = 11'd333;
      3: stateTransition = 11'd333;
      4: stateTransition = 11'd333;
      5: stateTransition = 11'd333;
      6: stateTransition = 11'd333;
      7: stateTransition = 11'd333;
      8: stateTransition = 11'd333;
      9: stateTransition = 11'd333;
      10: stateTransition = 11'd333;
      11: stateTransition = 11'd333;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd333;
      14: stateTransition = 11'd333;
      15: stateTransition = 11'd333;
      16: stateTransition = 11'd333;
      default: stateTransition = 11'bX;
    endcase
    334: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd334;
      2: stateTransition = 11'd334;
      3: stateTransition = 11'd334;
      4: stateTransition = 11'd334;
      5: stateTransition = 11'd334;
      6: stateTransition = 11'd334;
      7: stateTransition = 11'd334;
      8: stateTransition = 11'd334;
      9: stateTransition = 11'd334;
      10: stateTransition = 11'd334;
      11: stateTransition = 11'd334;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd334;
      14: stateTransition = 11'd334;
      15: stateTransition = 11'd334;
      16: stateTransition = 11'd334;
      default: stateTransition = 11'bX;
    endcase
    335: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd335;
      2: stateTransition = 11'd335;
      3: stateTransition = 11'd335;
      4: stateTransition = 11'd335;
      5: stateTransition = 11'd335;
      6: stateTransition = 11'd335;
      7: stateTransition = 11'd335;
      8: stateTransition = 11'd335;
      9: stateTransition = 11'd335;
      10: stateTransition = 11'd335;
      11: stateTransition = 11'd335;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd335;
      14: stateTransition = 11'd335;
      15: stateTransition = 11'd335;
      16: stateTransition = 11'd335;
      default: stateTransition = 11'bX;
    endcase
    336: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd336;
      2: stateTransition = 11'd336;
      3: stateTransition = 11'd336;
      4: stateTransition = 11'd336;
      5: stateTransition = 11'd336;
      6: stateTransition = 11'd336;
      7: stateTransition = 11'd336;
      8: stateTransition = 11'd336;
      9: stateTransition = 11'd336;
      10: stateTransition = 11'd336;
      11: stateTransition = 11'd336;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd336;
      14: stateTransition = 11'd336;
      15: stateTransition = 11'd336;
      16: stateTransition = 11'd336;
      default: stateTransition = 11'bX;
    endcase
    337: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd337;
      2: stateTransition = 11'd337;
      3: stateTransition = 11'd337;
      4: stateTransition = 11'd337;
      5: stateTransition = 11'd337;
      6: stateTransition = 11'd337;
      7: stateTransition = 11'd337;
      8: stateTransition = 11'd337;
      9: stateTransition = 11'd337;
      10: stateTransition = 11'd337;
      11: stateTransition = 11'd337;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd337;
      14: stateTransition = 11'd337;
      15: stateTransition = 11'd337;
      16: stateTransition = 11'd337;
      default: stateTransition = 11'bX;
    endcase
    338: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd338;
      2: stateTransition = 11'd338;
      3: stateTransition = 11'd338;
      4: stateTransition = 11'd338;
      5: stateTransition = 11'd338;
      6: stateTransition = 11'd338;
      7: stateTransition = 11'd338;
      8: stateTransition = 11'd338;
      9: stateTransition = 11'd338;
      10: stateTransition = 11'd338;
      11: stateTransition = 11'd338;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd338;
      14: stateTransition = 11'd338;
      15: stateTransition = 11'd338;
      16: stateTransition = 11'd338;
      default: stateTransition = 11'bX;
    endcase
    339: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd339;
      2: stateTransition = 11'd339;
      3: stateTransition = 11'd339;
      4: stateTransition = 11'd339;
      5: stateTransition = 11'd339;
      6: stateTransition = 11'd339;
      7: stateTransition = 11'd339;
      8: stateTransition = 11'd339;
      9: stateTransition = 11'd339;
      10: stateTransition = 11'd339;
      11: stateTransition = 11'd339;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd339;
      14: stateTransition = 11'd339;
      15: stateTransition = 11'd339;
      16: stateTransition = 11'd339;
      default: stateTransition = 11'bX;
    endcase
    340: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd340;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd340;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd340;
      8: stateTransition = 11'd340;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      default: stateTransition = 11'bX;
    endcase
    341: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd341;
      2: stateTransition = 11'd341;
      3: stateTransition = 11'd341;
      4: stateTransition = 11'd341;
      5: stateTransition = 11'd341;
      6: stateTransition = 11'd341;
      7: stateTransition = 11'd341;
      8: stateTransition = 11'd341;
      9: stateTransition = 11'd341;
      10: stateTransition = 11'd341;
      11: stateTransition = 11'd341;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd341;
      14: stateTransition = 11'd341;
      15: stateTransition = 11'd341;
      16: stateTransition = 11'd341;
      default: stateTransition = 11'bX;
    endcase
    342: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd342;
      2: stateTransition = 11'd342;
      3: stateTransition = 11'd342;
      4: stateTransition = 11'd342;
      5: stateTransition = 11'd342;
      6: stateTransition = 11'd342;
      7: stateTransition = 11'd342;
      8: stateTransition = 11'd342;
      9: stateTransition = 11'd342;
      10: stateTransition = 11'd342;
      11: stateTransition = 11'd342;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd342;
      14: stateTransition = 11'd342;
      15: stateTransition = 11'd342;
      16: stateTransition = 11'd342;
      default: stateTransition = 11'bX;
    endcase
    343: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd343;
      2: stateTransition = 11'd343;
      3: stateTransition = 11'd343;
      4: stateTransition = 11'd343;
      5: stateTransition = 11'd343;
      6: stateTransition = 11'd343;
      7: stateTransition = 11'd343;
      8: stateTransition = 11'd343;
      9: stateTransition = 11'd343;
      10: stateTransition = 11'd343;
      11: stateTransition = 11'd343;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd343;
      14: stateTransition = 11'd343;
      15: stateTransition = 11'd343;
      16: stateTransition = 11'd343;
      default: stateTransition = 11'bX;
    endcase
    344: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd344;
      2: stateTransition = 11'd344;
      3: stateTransition = 11'd344;
      4: stateTransition = 11'd344;
      5: stateTransition = 11'd344;
      6: stateTransition = 11'd344;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd344;
      10: stateTransition = 11'd344;
      11: stateTransition = 11'd344;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd344;
      14: stateTransition = 11'd344;
      15: stateTransition = 11'd344;
      16: stateTransition = 11'd344;
      default: stateTransition = 11'bX;
    endcase
    345: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd345;
      2: stateTransition = 11'd345;
      3: stateTransition = 11'd345;
      4: stateTransition = 11'd345;
      5: stateTransition = 11'd345;
      6: stateTransition = 11'd345;
      7: stateTransition = 11'd345;
      8: stateTransition = 11'd345;
      9: stateTransition = 11'd345;
      10: stateTransition = 11'd345;
      11: stateTransition = 11'd345;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd345;
      14: stateTransition = 11'd345;
      15: stateTransition = 11'd345;
      16: stateTransition = 11'd345;
      default: stateTransition = 11'bX;
    endcase
    346: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd346;
      2: stateTransition = 11'd346;
      3: stateTransition = 11'd346;
      4: stateTransition = 11'd346;
      5: stateTransition = 11'd346;
      6: stateTransition = 11'd346;
      7: stateTransition = 11'd346;
      8: stateTransition = 11'd346;
      9: stateTransition = 11'd346;
      10: stateTransition = 11'd346;
      11: stateTransition = 11'd346;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd346;
      14: stateTransition = 11'd346;
      15: stateTransition = 11'd346;
      16: stateTransition = 11'd346;
      default: stateTransition = 11'bX;
    endcase
    347: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd347;
      3: stateTransition = 11'd347;
      4: stateTransition = 11'd347;
      5: stateTransition = 11'd347;
      6: stateTransition = 11'd347;
      7: stateTransition = 11'd347;
      8: stateTransition = 11'd347;
      9: stateTransition = 11'd347;
      10: stateTransition = 11'd347;
      11: stateTransition = 11'd347;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd347;
      14: stateTransition = 11'd347;
      15: stateTransition = 11'd347;
      16: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    348: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd348;
      2: stateTransition = 11'd348;
      3: stateTransition = 11'd348;
      4: stateTransition = 11'd348;
      5: stateTransition = 11'd348;
      6: stateTransition = 11'd348;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd348;
      10: stateTransition = 11'd348;
      11: stateTransition = 11'd348;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd348;
      14: stateTransition = 11'd348;
      15: stateTransition = 11'd348;
      16: stateTransition = 11'd348;
      default: stateTransition = 11'bX;
    endcase
    349: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd349;
      2: stateTransition = 11'd349;
      3: stateTransition = 11'd349;
      4: stateTransition = 11'd349;
      5: stateTransition = 11'd349;
      6: stateTransition = 11'd349;
      7: stateTransition = 11'd349;
      8: stateTransition = 11'd349;
      9: stateTransition = 11'd349;
      10: stateTransition = 11'd349;
      11: stateTransition = 11'd349;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd349;
      14: stateTransition = 11'd349;
      15: stateTransition = 11'd349;
      16: stateTransition = 11'd349;
      default: stateTransition = 11'bX;
    endcase
    350: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd350;
      2: stateTransition = 11'd350;
      3: stateTransition = 11'd350;
      4: stateTransition = 11'd350;
      5: stateTransition = 11'd350;
      6: stateTransition = 11'd350;
      7: stateTransition = 11'd350;
      8: stateTransition = 11'd350;
      9: stateTransition = 11'd350;
      10: stateTransition = 11'd350;
      11: stateTransition = 11'd350;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd350;
      14: stateTransition = 11'd350;
      15: stateTransition = 11'd350;
      16: stateTransition = 11'd350;
      default: stateTransition = 11'bX;
    endcase
    351: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd351;
      2: stateTransition = 11'd351;
      3: stateTransition = 11'd351;
      4: stateTransition = 11'd351;
      5: stateTransition = 11'd351;
      6: stateTransition = 11'd351;
      7: stateTransition = 11'd351;
      8: stateTransition = 11'd351;
      9: stateTransition = 11'd351;
      10: stateTransition = 11'd351;
      11: stateTransition = 11'd351;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd351;
      14: stateTransition = 11'd351;
      15: stateTransition = 11'd351;
      16: stateTransition = 11'd351;
      default: stateTransition = 11'bX;
    endcase
    352: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd352;
      2: stateTransition = 11'd352;
      3: stateTransition = 11'd352;
      4: stateTransition = 11'd352;
      5: stateTransition = 11'd352;
      6: stateTransition = 11'd352;
      7: stateTransition = 11'd352;
      8: stateTransition = 11'd352;
      9: stateTransition = 11'd352;
      10: stateTransition = 11'd352;
      11: stateTransition = 11'd352;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd352;
      14: stateTransition = 11'd352;
      15: stateTransition = 11'd352;
      16: stateTransition = 11'd352;
      default: stateTransition = 11'bX;
    endcase
    353: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd353;
      2: stateTransition = 11'd353;
      3: stateTransition = 11'd353;
      4: stateTransition = 11'd353;
      5: stateTransition = 11'd353;
      6: stateTransition = 11'd353;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd353;
      9: stateTransition = 11'd353;
      10: stateTransition = 11'd353;
      11: stateTransition = 11'd353;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd353;
      14: stateTransition = 11'd353;
      15: stateTransition = 11'd353;
      16: stateTransition = 11'd353;
      default: stateTransition = 11'bX;
    endcase
    354: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd354;
      2: stateTransition = 11'd354;
      3: stateTransition = 11'd354;
      4: stateTransition = 11'd354;
      5: stateTransition = 11'd354;
      6: stateTransition = 11'd354;
      7: stateTransition = 11'd354;
      8: stateTransition = 11'd354;
      9: stateTransition = 11'd354;
      10: stateTransition = 11'd354;
      11: stateTransition = 11'd354;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd354;
      14: stateTransition = 11'd354;
      15: stateTransition = 11'd354;
      16: stateTransition = 11'd354;
      default: stateTransition = 11'bX;
    endcase
    355: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd355;
      2: stateTransition = 11'd355;
      3: stateTransition = 11'd355;
      4: stateTransition = 11'd355;
      5: stateTransition = 11'd355;
      6: stateTransition = 11'd355;
      7: stateTransition = 11'd355;
      8: stateTransition = 11'd355;
      9: stateTransition = 11'd355;
      10: stateTransition = 11'd355;
      11: stateTransition = 11'd355;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd355;
      14: stateTransition = 11'd355;
      15: stateTransition = 11'd355;
      16: stateTransition = 11'd355;
      default: stateTransition = 11'bX;
    endcase
    356: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd356;
      2: stateTransition = 11'd356;
      3: stateTransition = 11'd356;
      4: stateTransition = 11'd356;
      5: stateTransition = 11'd356;
      6: stateTransition = 11'd356;
      7: stateTransition = 11'd356;
      8: stateTransition = 11'd356;
      9: stateTransition = 11'd356;
      10: stateTransition = 11'd356;
      11: stateTransition = 11'd356;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd356;
      14: stateTransition = 11'd356;
      15: stateTransition = 11'd356;
      16: stateTransition = 11'd356;
      default: stateTransition = 11'bX;
    endcase
    357: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd357;
      2: stateTransition = 11'd357;
      3: stateTransition = 11'd357;
      4: stateTransition = 11'd357;
      5: stateTransition = 11'd357;
      6: stateTransition = 11'd357;
      7: stateTransition = 11'd357;
      8: stateTransition = 11'd357;
      9: stateTransition = 11'd357;
      10: stateTransition = 11'd357;
      11: stateTransition = 11'd357;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd357;
      14: stateTransition = 11'd357;
      15: stateTransition = 11'd357;
      16: stateTransition = 11'd357;
      default: stateTransition = 11'bX;
    endcase
    358: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    359: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd359;
      2: stateTransition = 11'd359;
      3: stateTransition = 11'd359;
      4: stateTransition = 11'd359;
      5: stateTransition = 11'd359;
      6: stateTransition = 11'd359;
      7: stateTransition = 11'd359;
      8: stateTransition = 11'd359;
      9: stateTransition = 11'd359;
      10: stateTransition = 11'd359;
      11: stateTransition = 11'd359;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd359;
      14: stateTransition = 11'd359;
      15: stateTransition = 11'd359;
      16: stateTransition = 11'd359;
      default: stateTransition = 11'bX;
    endcase
    360: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd360;
      2: stateTransition = 11'd360;
      3: stateTransition = 11'd360;
      4: stateTransition = 11'd360;
      5: stateTransition = 11'd360;
      6: stateTransition = 11'd360;
      7: stateTransition = 11'd360;
      8: stateTransition = 11'd360;
      9: stateTransition = 11'd360;
      10: stateTransition = 11'd360;
      11: stateTransition = 11'd360;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd360;
      14: stateTransition = 11'd360;
      15: stateTransition = 11'd360;
      16: stateTransition = 11'd360;
      default: stateTransition = 11'bX;
    endcase
    361: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd361;
      2: stateTransition = 11'd361;
      3: stateTransition = 11'd361;
      4: stateTransition = 11'd361;
      5: stateTransition = 11'd361;
      6: stateTransition = 11'd361;
      7: stateTransition = 11'd361;
      8: stateTransition = 11'd361;
      9: stateTransition = 11'd361;
      10: stateTransition = 11'd361;
      11: stateTransition = 11'd361;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd361;
      14: stateTransition = 11'd361;
      15: stateTransition = 11'd361;
      16: stateTransition = 11'd361;
      default: stateTransition = 11'bX;
    endcase
    362: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd362;
      2: stateTransition = 11'd362;
      3: stateTransition = 11'd362;
      4: stateTransition = 11'd362;
      5: stateTransition = 11'd362;
      6: stateTransition = 11'd362;
      7: stateTransition = 11'd362;
      8: stateTransition = 11'd362;
      9: stateTransition = 11'd362;
      10: stateTransition = 11'd362;
      11: stateTransition = 11'd362;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd362;
      14: stateTransition = 11'd362;
      15: stateTransition = 11'd362;
      16: stateTransition = 11'd362;
      default: stateTransition = 11'bX;
    endcase
    363: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd363;
      3: stateTransition = 11'd363;
      4: stateTransition = 11'd363;
      5: stateTransition = 11'd363;
      6: stateTransition = 11'd363;
      7: stateTransition = 11'd363;
      8: stateTransition = 11'd363;
      9: stateTransition = 11'd363;
      10: stateTransition = 11'd363;
      11: stateTransition = 11'd363;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd363;
      14: stateTransition = 11'd363;
      15: stateTransition = 11'd363;
      16: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    364: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd364;
      2: stateTransition = 11'd364;
      3: stateTransition = 11'd364;
      4: stateTransition = 11'd364;
      5: stateTransition = 11'd364;
      6: stateTransition = 11'd364;
      7: stateTransition = 11'd364;
      8: stateTransition = 11'd364;
      9: stateTransition = 11'd364;
      10: stateTransition = 11'd364;
      11: stateTransition = 11'd364;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd364;
      14: stateTransition = 11'd364;
      15: stateTransition = 11'd364;
      16: stateTransition = 11'd364;
      default: stateTransition = 11'bX;
    endcase
    365: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd365;
      2: stateTransition = 11'd365;
      3: stateTransition = 11'd365;
      4: stateTransition = 11'd365;
      5: stateTransition = 11'd365;
      6: stateTransition = 11'd365;
      7: stateTransition = 11'd365;
      8: stateTransition = 11'd365;
      9: stateTransition = 11'd365;
      10: stateTransition = 11'd365;
      11: stateTransition = 11'd365;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd365;
      14: stateTransition = 11'd365;
      15: stateTransition = 11'd365;
      16: stateTransition = 11'd365;
      default: stateTransition = 11'bX;
    endcase
    366: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd366;
      2: stateTransition = 11'd366;
      3: stateTransition = 11'd366;
      4: stateTransition = 11'd366;
      5: stateTransition = 11'd366;
      6: stateTransition = 11'd366;
      7: stateTransition = 11'd366;
      8: stateTransition = 11'd366;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd366;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd366;
      default: stateTransition = 11'bX;
    endcase
    367: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd367;
      2: stateTransition = 11'd367;
      3: stateTransition = 11'd367;
      4: stateTransition = 11'd367;
      5: stateTransition = 11'd367;
      6: stateTransition = 11'd367;
      7: stateTransition = 11'd367;
      8: stateTransition = 11'd367;
      9: stateTransition = 11'd367;
      10: stateTransition = 11'd367;
      11: stateTransition = 11'd367;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd367;
      14: stateTransition = 11'd367;
      15: stateTransition = 11'd367;
      16: stateTransition = 11'd367;
      default: stateTransition = 11'bX;
    endcase
    368: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd368;
      2: stateTransition = 11'd368;
      3: stateTransition = 11'd368;
      4: stateTransition = 11'd368;
      5: stateTransition = 11'd368;
      6: stateTransition = 11'd368;
      7: stateTransition = 11'd368;
      8: stateTransition = 11'd368;
      9: stateTransition = 11'd368;
      10: stateTransition = 11'd368;
      11: stateTransition = 11'd368;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd368;
      14: stateTransition = 11'd368;
      15: stateTransition = 11'd368;
      16: stateTransition = 11'd368;
      default: stateTransition = 11'bX;
    endcase
    369: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd369;
      5: stateTransition = 11'd369;
      6: stateTransition = 11'd369;
      7: stateTransition = 11'd369;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd369;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    370: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd370;
      2: stateTransition = 11'd370;
      3: stateTransition = 11'd370;
      4: stateTransition = 11'd370;
      5: stateTransition = 11'd370;
      6: stateTransition = 11'd370;
      7: stateTransition = 11'd370;
      8: stateTransition = 11'd370;
      9: stateTransition = 11'd370;
      10: stateTransition = 11'd370;
      11: stateTransition = 11'd370;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd370;
      14: stateTransition = 11'd370;
      15: stateTransition = 11'd370;
      16: stateTransition = 11'd370;
      default: stateTransition = 11'bX;
    endcase
    371: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd371;
      2: stateTransition = 11'd371;
      3: stateTransition = 11'd371;
      4: stateTransition = 11'd371;
      5: stateTransition = 11'd371;
      6: stateTransition = 11'd371;
      7: stateTransition = 11'd371;
      8: stateTransition = 11'd371;
      9: stateTransition = 11'd371;
      10: stateTransition = 11'd371;
      11: stateTransition = 11'd371;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd371;
      14: stateTransition = 11'd371;
      15: stateTransition = 11'd371;
      16: stateTransition = 11'd371;
      default: stateTransition = 11'bX;
    endcase
    372: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd372;
      2: stateTransition = 11'd372;
      3: stateTransition = 11'd372;
      4: stateTransition = 11'd372;
      5: stateTransition = 11'd372;
      6: stateTransition = 11'd372;
      7: stateTransition = 11'd372;
      8: stateTransition = 11'd372;
      9: stateTransition = 11'd372;
      10: stateTransition = 11'd372;
      11: stateTransition = 11'd372;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd372;
      14: stateTransition = 11'd372;
      15: stateTransition = 11'd372;
      16: stateTransition = 11'd372;
      default: stateTransition = 11'bX;
    endcase
    373: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd373;
      2: stateTransition = 11'd373;
      3: stateTransition = 11'd373;
      4: stateTransition = 11'd373;
      5: stateTransition = 11'd373;
      6: stateTransition = 11'd373;
      7: stateTransition = 11'd373;
      8: stateTransition = 11'd373;
      9: stateTransition = 11'd373;
      10: stateTransition = 11'd373;
      11: stateTransition = 11'd373;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd373;
      14: stateTransition = 11'd373;
      15: stateTransition = 11'd373;
      16: stateTransition = 11'd373;
      default: stateTransition = 11'bX;
    endcase
    374: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd374;
      2: stateTransition = 11'd374;
      3: stateTransition = 11'd374;
      4: stateTransition = 11'd374;
      5: stateTransition = 11'd374;
      6: stateTransition = 11'd374;
      7: stateTransition = 11'd374;
      8: stateTransition = 11'd374;
      9: stateTransition = 11'd374;
      10: stateTransition = 11'd374;
      11: stateTransition = 11'd374;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd374;
      14: stateTransition = 11'd374;
      15: stateTransition = 11'd374;
      16: stateTransition = 11'd374;
      default: stateTransition = 11'bX;
    endcase
    375: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd375;
      2: stateTransition = 11'd375;
      3: stateTransition = 11'd375;
      4: stateTransition = 11'd375;
      5: stateTransition = 11'd375;
      6: stateTransition = 11'd375;
      7: stateTransition = 11'd375;
      8: stateTransition = 11'd375;
      9: stateTransition = 11'd375;
      10: stateTransition = 11'd375;
      11: stateTransition = 11'd375;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd375;
      14: stateTransition = 11'd375;
      15: stateTransition = 11'd375;
      16: stateTransition = 11'd375;
      default: stateTransition = 11'bX;
    endcase
    376: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd376;
      2: stateTransition = 11'd376;
      3: stateTransition = 11'd376;
      4: stateTransition = 11'd376;
      5: stateTransition = 11'd376;
      6: stateTransition = 11'd376;
      7: stateTransition = 11'd376;
      8: stateTransition = 11'd376;
      9: stateTransition = 11'd376;
      10: stateTransition = 11'd376;
      11: stateTransition = 11'd376;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd376;
      14: stateTransition = 11'd376;
      15: stateTransition = 11'd376;
      16: stateTransition = 11'd376;
      default: stateTransition = 11'bX;
    endcase
    377: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd377;
      2: stateTransition = 11'd377;
      3: stateTransition = 11'd377;
      4: stateTransition = 11'd377;
      5: stateTransition = 11'd377;
      6: stateTransition = 11'd377;
      7: stateTransition = 11'd377;
      8: stateTransition = 11'd377;
      9: stateTransition = 11'd377;
      10: stateTransition = 11'd377;
      11: stateTransition = 11'd377;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd377;
      14: stateTransition = 11'd377;
      15: stateTransition = 11'd377;
      16: stateTransition = 11'd377;
      default: stateTransition = 11'bX;
    endcase
    378: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd378;
      2: stateTransition = 11'd378;
      3: stateTransition = 11'd378;
      4: stateTransition = 11'd378;
      5: stateTransition = 11'd378;
      6: stateTransition = 11'd378;
      7: stateTransition = 11'd378;
      8: stateTransition = 11'd378;
      9: stateTransition = 11'd378;
      10: stateTransition = 11'd378;
      11: stateTransition = 11'd378;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd378;
      14: stateTransition = 11'd378;
      15: stateTransition = 11'd378;
      16: stateTransition = 11'd378;
      default: stateTransition = 11'bX;
    endcase
    379: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd379;
      2: stateTransition = 11'd379;
      3: stateTransition = 11'd379;
      4: stateTransition = 11'd379;
      5: stateTransition = 11'd379;
      6: stateTransition = 11'd379;
      7: stateTransition = 11'd379;
      8: stateTransition = 11'd379;
      9: stateTransition = 11'd379;
      10: stateTransition = 11'd379;
      11: stateTransition = 11'd379;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd379;
      14: stateTransition = 11'd379;
      15: stateTransition = 11'd379;
      16: stateTransition = 11'd379;
      default: stateTransition = 11'bX;
    endcase
    380: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd380;
      2: stateTransition = 11'd380;
      3: stateTransition = 11'd380;
      4: stateTransition = 11'd380;
      5: stateTransition = 11'd380;
      6: stateTransition = 11'd380;
      7: stateTransition = 11'd380;
      8: stateTransition = 11'd380;
      9: stateTransition = 11'd380;
      10: stateTransition = 11'd380;
      11: stateTransition = 11'd380;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd380;
      14: stateTransition = 11'd380;
      15: stateTransition = 11'd380;
      16: stateTransition = 11'd380;
      default: stateTransition = 11'bX;
    endcase
    381: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd381;
      2: stateTransition = 11'd381;
      3: stateTransition = 11'd381;
      4: stateTransition = 11'd381;
      5: stateTransition = 11'd381;
      6: stateTransition = 11'd381;
      7: stateTransition = 11'd381;
      8: stateTransition = 11'd381;
      9: stateTransition = 11'd381;
      10: stateTransition = 11'd381;
      11: stateTransition = 11'd381;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd381;
      14: stateTransition = 11'd381;
      15: stateTransition = 11'd381;
      16: stateTransition = 11'd381;
      default: stateTransition = 11'bX;
    endcase
    382: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd382;
      2: stateTransition = 11'd382;
      3: stateTransition = 11'd382;
      4: stateTransition = 11'd382;
      5: stateTransition = 11'd382;
      6: stateTransition = 11'd382;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd382;
      9: stateTransition = 11'd382;
      10: stateTransition = 11'd382;
      11: stateTransition = 11'd382;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd382;
      14: stateTransition = 11'd382;
      15: stateTransition = 11'd382;
      16: stateTransition = 11'd382;
      default: stateTransition = 11'bX;
    endcase
    383: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd383;
      5: stateTransition = 11'd383;
      6: stateTransition = 11'd383;
      7: stateTransition = 11'd383;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd383;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    384: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd384;
      2: stateTransition = 11'd384;
      3: stateTransition = 11'd384;
      4: stateTransition = 11'd384;
      5: stateTransition = 11'd384;
      6: stateTransition = 11'd384;
      7: stateTransition = 11'd384;
      8: stateTransition = 11'd384;
      9: stateTransition = 11'd384;
      10: stateTransition = 11'd384;
      11: stateTransition = 11'd384;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd384;
      14: stateTransition = 11'd384;
      15: stateTransition = 11'd384;
      16: stateTransition = 11'd384;
      default: stateTransition = 11'bX;
    endcase
    385: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd385;
      2: stateTransition = 11'd385;
      3: stateTransition = 11'd385;
      4: stateTransition = 11'd385;
      5: stateTransition = 11'd385;
      6: stateTransition = 11'd385;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd385;
      9: stateTransition = 11'd385;
      10: stateTransition = 11'd385;
      11: stateTransition = 11'd385;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd385;
      14: stateTransition = 11'd385;
      15: stateTransition = 11'd385;
      16: stateTransition = 11'd385;
      default: stateTransition = 11'bX;
    endcase
    386: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd386;
      2: stateTransition = 11'd386;
      3: stateTransition = 11'd386;
      4: stateTransition = 11'd386;
      5: stateTransition = 11'd386;
      6: stateTransition = 11'd386;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd386;
      10: stateTransition = 11'd386;
      11: stateTransition = 11'd386;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd386;
      14: stateTransition = 11'd386;
      15: stateTransition = 11'd386;
      16: stateTransition = 11'd386;
      default: stateTransition = 11'bX;
    endcase
    387: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd387;
      2: stateTransition = 11'd387;
      3: stateTransition = 11'd387;
      4: stateTransition = 11'd387;
      5: stateTransition = 11'd387;
      6: stateTransition = 11'd387;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd387;
      10: stateTransition = 11'd387;
      11: stateTransition = 11'd387;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd387;
      14: stateTransition = 11'd387;
      15: stateTransition = 11'd387;
      16: stateTransition = 11'd387;
      default: stateTransition = 11'bX;
    endcase
    388: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd388;
      2: stateTransition = 11'd388;
      3: stateTransition = 11'd388;
      4: stateTransition = 11'd388;
      5: stateTransition = 11'd388;
      6: stateTransition = 11'd388;
      7: stateTransition = 11'd388;
      8: stateTransition = 11'd388;
      9: stateTransition = 11'd388;
      10: stateTransition = 11'd388;
      11: stateTransition = 11'd388;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd388;
      14: stateTransition = 11'd388;
      15: stateTransition = 11'd388;
      16: stateTransition = 11'd388;
      default: stateTransition = 11'bX;
    endcase
    389: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd389;
      2: stateTransition = 11'd389;
      3: stateTransition = 11'd389;
      4: stateTransition = 11'd389;
      5: stateTransition = 11'd389;
      6: stateTransition = 11'd389;
      7: stateTransition = 11'd389;
      8: stateTransition = 11'd389;
      9: stateTransition = 11'd389;
      10: stateTransition = 11'd389;
      11: stateTransition = 11'd389;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd389;
      14: stateTransition = 11'd389;
      15: stateTransition = 11'd389;
      16: stateTransition = 11'd389;
      default: stateTransition = 11'bX;
    endcase
    390: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd390;
      2: stateTransition = 11'd390;
      3: stateTransition = 11'd390;
      4: stateTransition = 11'd390;
      5: stateTransition = 11'd390;
      6: stateTransition = 11'd390;
      7: stateTransition = 11'd390;
      8: stateTransition = 11'd390;
      9: stateTransition = 11'd390;
      10: stateTransition = 11'd390;
      11: stateTransition = 11'd390;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd390;
      14: stateTransition = 11'd390;
      15: stateTransition = 11'd390;
      16: stateTransition = 11'd390;
      default: stateTransition = 11'bX;
    endcase
    391: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd391;
      2: stateTransition = 11'd391;
      3: stateTransition = 11'd391;
      4: stateTransition = 11'd391;
      5: stateTransition = 11'd391;
      6: stateTransition = 11'd391;
      7: stateTransition = 11'd391;
      8: stateTransition = 11'd391;
      9: stateTransition = 11'd391;
      10: stateTransition = 11'd391;
      11: stateTransition = 11'd391;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd391;
      14: stateTransition = 11'd391;
      15: stateTransition = 11'd391;
      16: stateTransition = 11'd391;
      default: stateTransition = 11'bX;
    endcase
    392: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd392;
      2: stateTransition = 11'd392;
      3: stateTransition = 11'd392;
      4: stateTransition = 11'd392;
      5: stateTransition = 11'd392;
      6: stateTransition = 11'd392;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd392;
      10: stateTransition = 11'd392;
      11: stateTransition = 11'd392;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd392;
      14: stateTransition = 11'd392;
      15: stateTransition = 11'd392;
      16: stateTransition = 11'd392;
      default: stateTransition = 11'bX;
    endcase
    393: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    394: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd394;
      2: stateTransition = 11'd394;
      3: stateTransition = 11'd394;
      4: stateTransition = 11'd394;
      5: stateTransition = 11'd394;
      6: stateTransition = 11'd394;
      7: stateTransition = 11'd394;
      8: stateTransition = 11'd394;
      9: stateTransition = 11'd394;
      10: stateTransition = 11'd394;
      11: stateTransition = 11'd394;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd394;
      14: stateTransition = 11'd394;
      15: stateTransition = 11'd394;
      16: stateTransition = 11'd394;
      default: stateTransition = 11'bX;
    endcase
    395: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd395;
      2: stateTransition = 11'd395;
      3: stateTransition = 11'd395;
      4: stateTransition = 11'd395;
      5: stateTransition = 11'd395;
      6: stateTransition = 11'd395;
      7: stateTransition = 11'd395;
      8: stateTransition = 11'd395;
      9: stateTransition = 11'd395;
      10: stateTransition = 11'd395;
      11: stateTransition = 11'd395;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd395;
      14: stateTransition = 11'd395;
      15: stateTransition = 11'd395;
      16: stateTransition = 11'd395;
      default: stateTransition = 11'bX;
    endcase
    396: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd396;
      2: stateTransition = 11'd396;
      3: stateTransition = 11'd396;
      4: stateTransition = 11'd396;
      5: stateTransition = 11'd396;
      6: stateTransition = 11'd396;
      7: stateTransition = 11'd396;
      8: stateTransition = 11'd396;
      9: stateTransition = 11'd396;
      10: stateTransition = 11'd396;
      11: stateTransition = 11'd396;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd396;
      14: stateTransition = 11'd396;
      15: stateTransition = 11'd396;
      16: stateTransition = 11'd396;
      default: stateTransition = 11'bX;
    endcase
    397: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd397;
      2: stateTransition = 11'd397;
      3: stateTransition = 11'd397;
      4: stateTransition = 11'd397;
      5: stateTransition = 11'd397;
      6: stateTransition = 11'd397;
      7: stateTransition = 11'd397;
      8: stateTransition = 11'd397;
      9: stateTransition = 11'd397;
      10: stateTransition = 11'd397;
      11: stateTransition = 11'd397;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd397;
      14: stateTransition = 11'd397;
      15: stateTransition = 11'd397;
      16: stateTransition = 11'd397;
      default: stateTransition = 11'bX;
    endcase
    398: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd398;
      2: stateTransition = 11'd398;
      3: stateTransition = 11'd398;
      4: stateTransition = 11'd398;
      5: stateTransition = 11'd398;
      6: stateTransition = 11'd398;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd398;
      9: stateTransition = 11'd398;
      10: stateTransition = 11'd398;
      11: stateTransition = 11'd398;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd398;
      14: stateTransition = 11'd398;
      15: stateTransition = 11'd398;
      16: stateTransition = 11'd398;
      default: stateTransition = 11'bX;
    endcase
    399: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd399;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd399;
      5: stateTransition = 11'd399;
      6: stateTransition = 11'd399;
      7: stateTransition = 11'd399;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd399;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    400: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd400;
      3: stateTransition = 11'd400;
      4: stateTransition = 11'd400;
      5: stateTransition = 11'd400;
      6: stateTransition = 11'd400;
      7: stateTransition = 11'd400;
      8: stateTransition = 11'd400;
      9: stateTransition = 11'd400;
      10: stateTransition = 11'd400;
      11: stateTransition = 11'd400;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd400;
      14: stateTransition = 11'd400;
      15: stateTransition = 11'd400;
      16: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    401: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd401;
      3: stateTransition = 11'd401;
      4: stateTransition = 11'd401;
      5: stateTransition = 11'd401;
      6: stateTransition = 11'd401;
      7: stateTransition = 11'd401;
      8: stateTransition = 11'd401;
      9: stateTransition = 11'd401;
      10: stateTransition = 11'd401;
      11: stateTransition = 11'd401;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd401;
      14: stateTransition = 11'd401;
      15: stateTransition = 11'd401;
      16: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    402: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd402;
      2: stateTransition = 11'd402;
      3: stateTransition = 11'd402;
      4: stateTransition = 11'd402;
      5: stateTransition = 11'd402;
      6: stateTransition = 11'd402;
      7: stateTransition = 11'd402;
      8: stateTransition = 11'd402;
      9: stateTransition = 11'd402;
      10: stateTransition = 11'd402;
      11: stateTransition = 11'd402;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd402;
      14: stateTransition = 11'd402;
      15: stateTransition = 11'd402;
      16: stateTransition = 11'd402;
      default: stateTransition = 11'bX;
    endcase
    403: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd403;
      2: stateTransition = 11'd403;
      3: stateTransition = 11'd403;
      4: stateTransition = 11'd403;
      5: stateTransition = 11'd403;
      6: stateTransition = 11'd403;
      7: stateTransition = 11'd403;
      8: stateTransition = 11'd403;
      9: stateTransition = 11'd403;
      10: stateTransition = 11'd403;
      11: stateTransition = 11'd403;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd403;
      14: stateTransition = 11'd403;
      15: stateTransition = 11'd403;
      16: stateTransition = 11'd403;
      default: stateTransition = 11'bX;
    endcase
    404: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd404;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd404;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd404;
      8: stateTransition = 11'd404;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      default: stateTransition = 11'bX;
    endcase
    405: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd405;
      2: stateTransition = 11'd405;
      3: stateTransition = 11'd405;
      4: stateTransition = 11'd405;
      5: stateTransition = 11'd405;
      6: stateTransition = 11'd405;
      7: stateTransition = 11'd405;
      8: stateTransition = 11'd405;
      9: stateTransition = 11'd405;
      10: stateTransition = 11'd405;
      11: stateTransition = 11'd405;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd405;
      14: stateTransition = 11'd405;
      15: stateTransition = 11'd405;
      16: stateTransition = 11'd405;
      default: stateTransition = 11'bX;
    endcase
    406: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd406;
      2: stateTransition = 11'd406;
      3: stateTransition = 11'd406;
      4: stateTransition = 11'd406;
      5: stateTransition = 11'd406;
      6: stateTransition = 11'd406;
      7: stateTransition = 11'd406;
      8: stateTransition = 11'd406;
      9: stateTransition = 11'd406;
      10: stateTransition = 11'd406;
      11: stateTransition = 11'd406;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd406;
      14: stateTransition = 11'd406;
      15: stateTransition = 11'd406;
      16: stateTransition = 11'd406;
      default: stateTransition = 11'bX;
    endcase
    407: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd407;
      2: stateTransition = 11'd407;
      3: stateTransition = 11'd407;
      4: stateTransition = 11'd407;
      5: stateTransition = 11'd407;
      6: stateTransition = 11'd407;
      7: stateTransition = 11'd407;
      8: stateTransition = 11'd407;
      9: stateTransition = 11'd407;
      10: stateTransition = 11'd407;
      11: stateTransition = 11'd407;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd407;
      14: stateTransition = 11'd407;
      15: stateTransition = 11'd407;
      16: stateTransition = 11'd407;
      default: stateTransition = 11'bX;
    endcase
    408: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd408;
      2: stateTransition = 11'd408;
      3: stateTransition = 11'd408;
      4: stateTransition = 11'd408;
      5: stateTransition = 11'd408;
      6: stateTransition = 11'd408;
      7: stateTransition = 11'd408;
      8: stateTransition = 11'd408;
      9: stateTransition = 11'd408;
      10: stateTransition = 11'd408;
      11: stateTransition = 11'd408;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd408;
      14: stateTransition = 11'd408;
      15: stateTransition = 11'd408;
      16: stateTransition = 11'd408;
      default: stateTransition = 11'bX;
    endcase
    409: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd409;
      2: stateTransition = 11'd409;
      3: stateTransition = 11'd409;
      4: stateTransition = 11'd409;
      5: stateTransition = 11'd409;
      6: stateTransition = 11'd409;
      7: stateTransition = 11'd409;
      8: stateTransition = 11'd409;
      9: stateTransition = 11'd409;
      10: stateTransition = 11'd409;
      11: stateTransition = 11'd409;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd409;
      14: stateTransition = 11'd409;
      15: stateTransition = 11'd409;
      16: stateTransition = 11'd409;
      default: stateTransition = 11'bX;
    endcase
    410: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd410;
      2: stateTransition = 11'd410;
      3: stateTransition = 11'd410;
      4: stateTransition = 11'd410;
      5: stateTransition = 11'd410;
      6: stateTransition = 11'd410;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd410;
      9: stateTransition = 11'd410;
      10: stateTransition = 11'd410;
      11: stateTransition = 11'd410;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd410;
      14: stateTransition = 11'd410;
      15: stateTransition = 11'd410;
      16: stateTransition = 11'd410;
      default: stateTransition = 11'bX;
    endcase
    411: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd411;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd411;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    412: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd412;
      2: stateTransition = 11'd412;
      3: stateTransition = 11'd412;
      4: stateTransition = 11'd412;
      5: stateTransition = 11'd412;
      6: stateTransition = 11'd412;
      7: stateTransition = 11'd412;
      8: stateTransition = 11'd412;
      9: stateTransition = 11'd412;
      10: stateTransition = 11'd412;
      11: stateTransition = 11'd412;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd412;
      14: stateTransition = 11'd412;
      15: stateTransition = 11'd412;
      16: stateTransition = 11'd412;
      default: stateTransition = 11'bX;
    endcase
    413: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd413;
      2: stateTransition = 11'd413;
      3: stateTransition = 11'd413;
      4: stateTransition = 11'd413;
      5: stateTransition = 11'd413;
      6: stateTransition = 11'd413;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd413;
      9: stateTransition = 11'd413;
      10: stateTransition = 11'd413;
      11: stateTransition = 11'd413;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd413;
      14: stateTransition = 11'd413;
      15: stateTransition = 11'd413;
      16: stateTransition = 11'd413;
      default: stateTransition = 11'bX;
    endcase
    414: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd414;
      2: stateTransition = 11'd414;
      3: stateTransition = 11'd414;
      4: stateTransition = 11'd414;
      5: stateTransition = 11'd414;
      6: stateTransition = 11'd414;
      7: stateTransition = 11'd414;
      8: stateTransition = 11'd414;
      9: stateTransition = 11'd414;
      10: stateTransition = 11'd414;
      11: stateTransition = 11'd414;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd414;
      14: stateTransition = 11'd414;
      15: stateTransition = 11'd414;
      16: stateTransition = 11'd414;
      default: stateTransition = 11'bX;
    endcase
    415: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd415;
      2: stateTransition = 11'd415;
      3: stateTransition = 11'd415;
      4: stateTransition = 11'd415;
      5: stateTransition = 11'd415;
      6: stateTransition = 11'd415;
      7: stateTransition = 11'd415;
      8: stateTransition = 11'd415;
      9: stateTransition = 11'd415;
      10: stateTransition = 11'd415;
      11: stateTransition = 11'd415;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd415;
      14: stateTransition = 11'd415;
      15: stateTransition = 11'd415;
      16: stateTransition = 11'd415;
      default: stateTransition = 11'bX;
    endcase
    416: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd416;
      2: stateTransition = 11'd416;
      3: stateTransition = 11'd416;
      4: stateTransition = 11'd416;
      5: stateTransition = 11'd416;
      6: stateTransition = 11'd416;
      7: stateTransition = 11'd416;
      8: stateTransition = 11'd416;
      9: stateTransition = 11'd416;
      10: stateTransition = 11'd416;
      11: stateTransition = 11'd416;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd416;
      14: stateTransition = 11'd416;
      15: stateTransition = 11'd416;
      16: stateTransition = 11'd416;
      default: stateTransition = 11'bX;
    endcase
    417: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd417;
      2: stateTransition = 11'd417;
      3: stateTransition = 11'd417;
      4: stateTransition = 11'd417;
      5: stateTransition = 11'd417;
      6: stateTransition = 11'd417;
      7: stateTransition = 11'd417;
      8: stateTransition = 11'd417;
      9: stateTransition = 11'd417;
      10: stateTransition = 11'd417;
      11: stateTransition = 11'd417;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd417;
      14: stateTransition = 11'd417;
      15: stateTransition = 11'd417;
      16: stateTransition = 11'd417;
      default: stateTransition = 11'bX;
    endcase
    418: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd418;
      2: stateTransition = 11'd418;
      3: stateTransition = 11'd418;
      4: stateTransition = 11'd418;
      5: stateTransition = 11'd418;
      6: stateTransition = 11'd418;
      7: stateTransition = 11'd418;
      8: stateTransition = 11'd418;
      9: stateTransition = 11'd418;
      10: stateTransition = 11'd418;
      11: stateTransition = 11'd418;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd418;
      14: stateTransition = 11'd418;
      15: stateTransition = 11'd418;
      16: stateTransition = 11'd418;
      default: stateTransition = 11'bX;
    endcase
    419: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd419;
      2: stateTransition = 11'd419;
      3: stateTransition = 11'd419;
      4: stateTransition = 11'd419;
      5: stateTransition = 11'd419;
      6: stateTransition = 11'd419;
      7: stateTransition = 11'd419;
      8: stateTransition = 11'd419;
      9: stateTransition = 11'd419;
      10: stateTransition = 11'd419;
      11: stateTransition = 11'd419;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd419;
      14: stateTransition = 11'd419;
      15: stateTransition = 11'd419;
      16: stateTransition = 11'd419;
      default: stateTransition = 11'bX;
    endcase
    420: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd420;
      2: stateTransition = 11'd420;
      3: stateTransition = 11'd420;
      4: stateTransition = 11'd420;
      5: stateTransition = 11'd420;
      6: stateTransition = 11'd420;
      7: stateTransition = 11'd420;
      8: stateTransition = 11'd420;
      9: stateTransition = 11'd420;
      10: stateTransition = 11'd420;
      11: stateTransition = 11'd420;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd420;
      14: stateTransition = 11'd420;
      15: stateTransition = 11'd420;
      16: stateTransition = 11'd420;
      default: stateTransition = 11'bX;
    endcase
    421: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd421;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd421;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd421;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd421;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd421;
      16: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    422: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd422;
      2: stateTransition = 11'd422;
      3: stateTransition = 11'd422;
      4: stateTransition = 11'd422;
      5: stateTransition = 11'd422;
      6: stateTransition = 11'd422;
      7: stateTransition = 11'd422;
      8: stateTransition = 11'd422;
      9: stateTransition = 11'd422;
      10: stateTransition = 11'd422;
      11: stateTransition = 11'd422;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd422;
      14: stateTransition = 11'd422;
      15: stateTransition = 11'd422;
      16: stateTransition = 11'd422;
      default: stateTransition = 11'bX;
    endcase
    423: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd423;
      2: stateTransition = 11'd423;
      3: stateTransition = 11'd423;
      4: stateTransition = 11'd423;
      5: stateTransition = 11'd423;
      6: stateTransition = 11'd423;
      7: stateTransition = 11'd423;
      8: stateTransition = 11'd423;
      9: stateTransition = 11'd423;
      10: stateTransition = 11'd423;
      11: stateTransition = 11'd423;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd423;
      14: stateTransition = 11'd423;
      15: stateTransition = 11'd423;
      16: stateTransition = 11'd423;
      default: stateTransition = 11'bX;
    endcase
    424: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd424;
      2: stateTransition = 11'd424;
      3: stateTransition = 11'd424;
      4: stateTransition = 11'd424;
      5: stateTransition = 11'd424;
      6: stateTransition = 11'd424;
      7: stateTransition = 11'd424;
      8: stateTransition = 11'd424;
      9: stateTransition = 11'd424;
      10: stateTransition = 11'd424;
      11: stateTransition = 11'd424;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd424;
      14: stateTransition = 11'd424;
      15: stateTransition = 11'd424;
      16: stateTransition = 11'd424;
      default: stateTransition = 11'bX;
    endcase
    425: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd425;
      2: stateTransition = 11'd425;
      3: stateTransition = 11'd425;
      4: stateTransition = 11'd425;
      5: stateTransition = 11'd425;
      6: stateTransition = 11'd425;
      7: stateTransition = 11'd425;
      8: stateTransition = 11'd425;
      9: stateTransition = 11'd425;
      10: stateTransition = 11'd425;
      11: stateTransition = 11'd425;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd425;
      14: stateTransition = 11'd425;
      15: stateTransition = 11'd425;
      16: stateTransition = 11'd425;
      default: stateTransition = 11'bX;
    endcase
    426: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd426;
      2: stateTransition = 11'd426;
      3: stateTransition = 11'd426;
      4: stateTransition = 11'd426;
      5: stateTransition = 11'd426;
      6: stateTransition = 11'd426;
      7: stateTransition = 11'd426;
      8: stateTransition = 11'd426;
      9: stateTransition = 11'd426;
      10: stateTransition = 11'd426;
      11: stateTransition = 11'd426;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd426;
      14: stateTransition = 11'd426;
      15: stateTransition = 11'd426;
      16: stateTransition = 11'd426;
      default: stateTransition = 11'bX;
    endcase
    427: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd427;
      2: stateTransition = 11'd427;
      3: stateTransition = 11'd427;
      4: stateTransition = 11'd427;
      5: stateTransition = 11'd427;
      6: stateTransition = 11'd427;
      7: stateTransition = 11'd427;
      8: stateTransition = 11'd427;
      9: stateTransition = 11'd427;
      10: stateTransition = 11'd427;
      11: stateTransition = 11'd427;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd427;
      14: stateTransition = 11'd427;
      15: stateTransition = 11'd427;
      16: stateTransition = 11'd427;
      default: stateTransition = 11'bX;
    endcase
    428: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd428;
      2: stateTransition = 11'd428;
      3: stateTransition = 11'd428;
      4: stateTransition = 11'd428;
      5: stateTransition = 11'd428;
      6: stateTransition = 11'd428;
      7: stateTransition = 11'd428;
      8: stateTransition = 11'd428;
      9: stateTransition = 11'd428;
      10: stateTransition = 11'd428;
      11: stateTransition = 11'd428;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd428;
      14: stateTransition = 11'd428;
      15: stateTransition = 11'd428;
      16: stateTransition = 11'd428;
      default: stateTransition = 11'bX;
    endcase
    429: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd429;
      2: stateTransition = 11'd429;
      3: stateTransition = 11'd429;
      4: stateTransition = 11'd429;
      5: stateTransition = 11'd429;
      6: stateTransition = 11'd429;
      7: stateTransition = 11'd429;
      8: stateTransition = 11'd429;
      9: stateTransition = 11'd429;
      10: stateTransition = 11'd429;
      11: stateTransition = 11'd429;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd429;
      14: stateTransition = 11'd429;
      15: stateTransition = 11'd429;
      16: stateTransition = 11'd429;
      default: stateTransition = 11'bX;
    endcase
    430: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd430;
      2: stateTransition = 11'd430;
      3: stateTransition = 11'd430;
      4: stateTransition = 11'd430;
      5: stateTransition = 11'd430;
      6: stateTransition = 11'd430;
      7: stateTransition = 11'd430;
      8: stateTransition = 11'd430;
      9: stateTransition = 11'd430;
      10: stateTransition = 11'd430;
      11: stateTransition = 11'd430;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd430;
      14: stateTransition = 11'd430;
      15: stateTransition = 11'd430;
      16: stateTransition = 11'd430;
      default: stateTransition = 11'bX;
    endcase
    431: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd431;
      2: stateTransition = 11'd431;
      3: stateTransition = 11'd431;
      4: stateTransition = 11'd431;
      5: stateTransition = 11'd431;
      6: stateTransition = 11'd431;
      7: stateTransition = 11'd431;
      8: stateTransition = 11'd431;
      9: stateTransition = 11'd431;
      10: stateTransition = 11'd431;
      11: stateTransition = 11'd431;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd431;
      14: stateTransition = 11'd431;
      15: stateTransition = 11'd431;
      16: stateTransition = 11'd431;
      default: stateTransition = 11'bX;
    endcase
    432: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd432;
      2: stateTransition = 11'd432;
      3: stateTransition = 11'd432;
      4: stateTransition = 11'd432;
      5: stateTransition = 11'd432;
      6: stateTransition = 11'd432;
      7: stateTransition = 11'd432;
      8: stateTransition = 11'd432;
      9: stateTransition = 11'd432;
      10: stateTransition = 11'd432;
      11: stateTransition = 11'd432;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd432;
      14: stateTransition = 11'd432;
      15: stateTransition = 11'd432;
      16: stateTransition = 11'd432;
      default: stateTransition = 11'bX;
    endcase
    433: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd433;
      2: stateTransition = 11'd433;
      3: stateTransition = 11'd433;
      4: stateTransition = 11'd433;
      5: stateTransition = 11'd433;
      6: stateTransition = 11'd433;
      7: stateTransition = 11'd433;
      8: stateTransition = 11'd433;
      9: stateTransition = 11'd433;
      10: stateTransition = 11'd433;
      11: stateTransition = 11'd433;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd433;
      14: stateTransition = 11'd433;
      15: stateTransition = 11'd433;
      16: stateTransition = 11'd433;
      default: stateTransition = 11'bX;
    endcase
    434: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd434;
      2: stateTransition = 11'd434;
      3: stateTransition = 11'd434;
      4: stateTransition = 11'd434;
      5: stateTransition = 11'd434;
      6: stateTransition = 11'd434;
      7: stateTransition = 11'd434;
      8: stateTransition = 11'd434;
      9: stateTransition = 11'd434;
      10: stateTransition = 11'd434;
      11: stateTransition = 11'd434;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd434;
      14: stateTransition = 11'd434;
      15: stateTransition = 11'd434;
      16: stateTransition = 11'd434;
      default: stateTransition = 11'bX;
    endcase
    435: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd435;
      2: stateTransition = 11'd435;
      3: stateTransition = 11'd435;
      4: stateTransition = 11'd435;
      5: stateTransition = 11'd435;
      6: stateTransition = 11'd435;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd435;
      9: stateTransition = 11'd435;
      10: stateTransition = 11'd435;
      11: stateTransition = 11'd435;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd435;
      14: stateTransition = 11'd435;
      15: stateTransition = 11'd435;
      16: stateTransition = 11'd435;
      default: stateTransition = 11'bX;
    endcase
    436: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd436;
      5: stateTransition = 11'd436;
      6: stateTransition = 11'd436;
      7: stateTransition = 11'd436;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd436;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    437: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd437;
      2: stateTransition = 11'd437;
      3: stateTransition = 11'd437;
      4: stateTransition = 11'd437;
      5: stateTransition = 11'd437;
      6: stateTransition = 11'd437;
      7: stateTransition = 11'd437;
      8: stateTransition = 11'd437;
      9: stateTransition = 11'd437;
      10: stateTransition = 11'd437;
      11: stateTransition = 11'd437;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd437;
      14: stateTransition = 11'd437;
      15: stateTransition = 11'd437;
      16: stateTransition = 11'd437;
      default: stateTransition = 11'bX;
    endcase
    438: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd438;
      2: stateTransition = 11'd438;
      3: stateTransition = 11'd438;
      4: stateTransition = 11'd438;
      5: stateTransition = 11'd438;
      6: stateTransition = 11'd438;
      7: stateTransition = 11'd438;
      8: stateTransition = 11'd438;
      9: stateTransition = 11'd438;
      10: stateTransition = 11'd438;
      11: stateTransition = 11'd438;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd438;
      14: stateTransition = 11'd438;
      15: stateTransition = 11'd438;
      16: stateTransition = 11'd438;
      default: stateTransition = 11'bX;
    endcase
    439: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd439;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd439;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd439;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd439;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd439;
      16: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    440: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd440;
      2: stateTransition = 11'd440;
      3: stateTransition = 11'd440;
      4: stateTransition = 11'd440;
      5: stateTransition = 11'd440;
      6: stateTransition = 11'd440;
      7: stateTransition = 11'd440;
      8: stateTransition = 11'd440;
      9: stateTransition = 11'd440;
      10: stateTransition = 11'd440;
      11: stateTransition = 11'd440;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd440;
      14: stateTransition = 11'd440;
      15: stateTransition = 11'd440;
      16: stateTransition = 11'd440;
      default: stateTransition = 11'bX;
    endcase
    441: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd441;
      2: stateTransition = 11'd441;
      3: stateTransition = 11'd441;
      4: stateTransition = 11'd441;
      5: stateTransition = 11'd441;
      6: stateTransition = 11'd441;
      7: stateTransition = 11'd441;
      8: stateTransition = 11'd441;
      9: stateTransition = 11'd441;
      10: stateTransition = 11'd441;
      11: stateTransition = 11'd441;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd441;
      14: stateTransition = 11'd441;
      15: stateTransition = 11'd441;
      16: stateTransition = 11'd441;
      default: stateTransition = 11'bX;
    endcase
    442: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd442;
      2: stateTransition = 11'd442;
      3: stateTransition = 11'd442;
      4: stateTransition = 11'd442;
      5: stateTransition = 11'd442;
      6: stateTransition = 11'd442;
      7: stateTransition = 11'd442;
      8: stateTransition = 11'd442;
      9: stateTransition = 11'd442;
      10: stateTransition = 11'd442;
      11: stateTransition = 11'd442;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd442;
      14: stateTransition = 11'd442;
      15: stateTransition = 11'd442;
      16: stateTransition = 11'd442;
      default: stateTransition = 11'bX;
    endcase
    443: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd443;
      2: stateTransition = 11'd443;
      3: stateTransition = 11'd443;
      4: stateTransition = 11'd443;
      5: stateTransition = 11'd443;
      6: stateTransition = 11'd443;
      7: stateTransition = 11'd443;
      8: stateTransition = 11'd443;
      9: stateTransition = 11'd443;
      10: stateTransition = 11'd443;
      11: stateTransition = 11'd443;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd443;
      14: stateTransition = 11'd443;
      15: stateTransition = 11'd443;
      16: stateTransition = 11'd443;
      default: stateTransition = 11'bX;
    endcase
    444: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd444;
      2: stateTransition = 11'd444;
      3: stateTransition = 11'd444;
      4: stateTransition = 11'd444;
      5: stateTransition = 11'd444;
      6: stateTransition = 11'd444;
      7: stateTransition = 11'd444;
      8: stateTransition = 11'd444;
      9: stateTransition = 11'd444;
      10: stateTransition = 11'd444;
      11: stateTransition = 11'd444;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd444;
      14: stateTransition = 11'd444;
      15: stateTransition = 11'd444;
      16: stateTransition = 11'd444;
      default: stateTransition = 11'bX;
    endcase
    445: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd445;
      2: stateTransition = 11'd445;
      3: stateTransition = 11'd445;
      4: stateTransition = 11'd445;
      5: stateTransition = 11'd445;
      6: stateTransition = 11'd445;
      7: stateTransition = 11'd445;
      8: stateTransition = 11'd445;
      9: stateTransition = 11'd445;
      10: stateTransition = 11'd445;
      11: stateTransition = 11'd445;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd445;
      14: stateTransition = 11'd445;
      15: stateTransition = 11'd445;
      16: stateTransition = 11'd445;
      default: stateTransition = 11'bX;
    endcase
    446: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd446;
      2: stateTransition = 11'd446;
      3: stateTransition = 11'd446;
      4: stateTransition = 11'd446;
      5: stateTransition = 11'd446;
      6: stateTransition = 11'd446;
      7: stateTransition = 11'd446;
      8: stateTransition = 11'd446;
      9: stateTransition = 11'd446;
      10: stateTransition = 11'd446;
      11: stateTransition = 11'd446;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd446;
      14: stateTransition = 11'd446;
      15: stateTransition = 11'd446;
      16: stateTransition = 11'd446;
      default: stateTransition = 11'bX;
    endcase
    447: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd447;
      2: stateTransition = 11'd447;
      3: stateTransition = 11'd447;
      4: stateTransition = 11'd447;
      5: stateTransition = 11'd447;
      6: stateTransition = 11'd447;
      7: stateTransition = 11'd447;
      8: stateTransition = 11'd447;
      9: stateTransition = 11'd447;
      10: stateTransition = 11'd447;
      11: stateTransition = 11'd447;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd447;
      14: stateTransition = 11'd447;
      15: stateTransition = 11'd447;
      16: stateTransition = 11'd447;
      default: stateTransition = 11'bX;
    endcase
    448: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd448;
      2: stateTransition = 11'd448;
      3: stateTransition = 11'd448;
      4: stateTransition = 11'd448;
      5: stateTransition = 11'd448;
      6: stateTransition = 11'd448;
      7: stateTransition = 11'd448;
      8: stateTransition = 11'd448;
      9: stateTransition = 11'd448;
      10: stateTransition = 11'd448;
      11: stateTransition = 11'd448;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd448;
      14: stateTransition = 11'd448;
      15: stateTransition = 11'd448;
      16: stateTransition = 11'd448;
      default: stateTransition = 11'bX;
    endcase
    449: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd449;
      2: stateTransition = 11'd449;
      3: stateTransition = 11'd449;
      4: stateTransition = 11'd449;
      5: stateTransition = 11'd449;
      6: stateTransition = 11'd449;
      7: stateTransition = 11'd449;
      8: stateTransition = 11'd449;
      9: stateTransition = 11'd449;
      10: stateTransition = 11'd449;
      11: stateTransition = 11'd449;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd449;
      14: stateTransition = 11'd449;
      15: stateTransition = 11'd449;
      16: stateTransition = 11'd449;
      default: stateTransition = 11'bX;
    endcase
    450: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd450;
      2: stateTransition = 11'd450;
      3: stateTransition = 11'd450;
      4: stateTransition = 11'd450;
      5: stateTransition = 11'd450;
      6: stateTransition = 11'd450;
      7: stateTransition = 11'd450;
      8: stateTransition = 11'd450;
      9: stateTransition = 11'd450;
      10: stateTransition = 11'd450;
      11: stateTransition = 11'd450;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd450;
      14: stateTransition = 11'd450;
      15: stateTransition = 11'd450;
      16: stateTransition = 11'd450;
      default: stateTransition = 11'bX;
    endcase
    451: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd451;
      2: stateTransition = 11'd451;
      3: stateTransition = 11'd451;
      4: stateTransition = 11'd451;
      5: stateTransition = 11'd451;
      6: stateTransition = 11'd451;
      7: stateTransition = 11'd451;
      8: stateTransition = 11'd451;
      9: stateTransition = 11'd451;
      10: stateTransition = 11'd451;
      11: stateTransition = 11'd451;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd451;
      14: stateTransition = 11'd451;
      15: stateTransition = 11'd451;
      16: stateTransition = 11'd451;
      default: stateTransition = 11'bX;
    endcase
    452: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd452;
      2: stateTransition = 11'd452;
      3: stateTransition = 11'd452;
      4: stateTransition = 11'd452;
      5: stateTransition = 11'd452;
      6: stateTransition = 11'd452;
      7: stateTransition = 11'd452;
      8: stateTransition = 11'd452;
      9: stateTransition = 11'd452;
      10: stateTransition = 11'd452;
      11: stateTransition = 11'd452;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd452;
      14: stateTransition = 11'd452;
      15: stateTransition = 11'd452;
      16: stateTransition = 11'd452;
      default: stateTransition = 11'bX;
    endcase
    453: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd453;
      2: stateTransition = 11'd453;
      3: stateTransition = 11'd453;
      4: stateTransition = 11'd453;
      5: stateTransition = 11'd453;
      6: stateTransition = 11'd453;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd453;
      9: stateTransition = 11'd453;
      10: stateTransition = 11'd453;
      11: stateTransition = 11'd453;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd453;
      14: stateTransition = 11'd453;
      15: stateTransition = 11'd453;
      16: stateTransition = 11'd453;
      default: stateTransition = 11'bX;
    endcase
    454: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd454;
      2: stateTransition = 11'd454;
      3: stateTransition = 11'd454;
      4: stateTransition = 11'd454;
      5: stateTransition = 11'd454;
      6: stateTransition = 11'd454;
      7: stateTransition = 11'd454;
      8: stateTransition = 11'd454;
      9: stateTransition = 11'd454;
      10: stateTransition = 11'd454;
      11: stateTransition = 11'd454;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd454;
      14: stateTransition = 11'd454;
      15: stateTransition = 11'd454;
      16: stateTransition = 11'd454;
      default: stateTransition = 11'bX;
    endcase
    455: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd455;
      5: stateTransition = 11'd455;
      6: stateTransition = 11'd455;
      7: stateTransition = 11'd455;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd455;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    456: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd456;
      2: stateTransition = 11'd456;
      3: stateTransition = 11'd456;
      4: stateTransition = 11'd456;
      5: stateTransition = 11'd456;
      6: stateTransition = 11'd456;
      7: stateTransition = 11'd456;
      8: stateTransition = 11'd456;
      9: stateTransition = 11'd456;
      10: stateTransition = 11'd456;
      11: stateTransition = 11'd456;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd456;
      14: stateTransition = 11'd456;
      15: stateTransition = 11'd456;
      16: stateTransition = 11'd456;
      default: stateTransition = 11'bX;
    endcase
    457: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd457;
      2: stateTransition = 11'd457;
      3: stateTransition = 11'd457;
      4: stateTransition = 11'd457;
      5: stateTransition = 11'd457;
      6: stateTransition = 11'd457;
      7: stateTransition = 11'd457;
      8: stateTransition = 11'd457;
      9: stateTransition = 11'd457;
      10: stateTransition = 11'd457;
      11: stateTransition = 11'd457;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd457;
      14: stateTransition = 11'd457;
      15: stateTransition = 11'd457;
      16: stateTransition = 11'd457;
      default: stateTransition = 11'bX;
    endcase
    458: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd458;
      2: stateTransition = 11'd458;
      3: stateTransition = 11'd458;
      4: stateTransition = 11'd458;
      5: stateTransition = 11'd458;
      6: stateTransition = 11'd458;
      7: stateTransition = 11'd458;
      8: stateTransition = 11'd458;
      9: stateTransition = 11'd458;
      10: stateTransition = 11'd458;
      11: stateTransition = 11'd458;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd458;
      14: stateTransition = 11'd458;
      15: stateTransition = 11'd458;
      16: stateTransition = 11'd458;
      default: stateTransition = 11'bX;
    endcase
    459: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd459;
      2: stateTransition = 11'd459;
      3: stateTransition = 11'd459;
      4: stateTransition = 11'd459;
      5: stateTransition = 11'd459;
      6: stateTransition = 11'd459;
      7: stateTransition = 11'd459;
      8: stateTransition = 11'd459;
      9: stateTransition = 11'd459;
      10: stateTransition = 11'd459;
      11: stateTransition = 11'd459;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd459;
      14: stateTransition = 11'd459;
      15: stateTransition = 11'd459;
      16: stateTransition = 11'd459;
      default: stateTransition = 11'bX;
    endcase
    460: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd460;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd460;
      10: stateTransition = 11'd460;
      11: stateTransition = 11'd460;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd460;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd460;
      16: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    461: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd461;
      2: stateTransition = 11'd461;
      3: stateTransition = 11'd461;
      4: stateTransition = 11'd461;
      5: stateTransition = 11'd461;
      6: stateTransition = 11'd461;
      7: stateTransition = 11'd461;
      8: stateTransition = 11'd461;
      9: stateTransition = 11'd461;
      10: stateTransition = 11'd461;
      11: stateTransition = 11'd461;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd461;
      14: stateTransition = 11'd461;
      15: stateTransition = 11'd461;
      16: stateTransition = 11'd461;
      default: stateTransition = 11'bX;
    endcase
    462: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd462;
      2: stateTransition = 11'd462;
      3: stateTransition = 11'd462;
      4: stateTransition = 11'd462;
      5: stateTransition = 11'd462;
      6: stateTransition = 11'd462;
      7: stateTransition = 11'd462;
      8: stateTransition = 11'd462;
      9: stateTransition = 11'd462;
      10: stateTransition = 11'd462;
      11: stateTransition = 11'd462;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd462;
      14: stateTransition = 11'd462;
      15: stateTransition = 11'd462;
      16: stateTransition = 11'd462;
      default: stateTransition = 11'bX;
    endcase
    463: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd463;
      2: stateTransition = 11'd463;
      3: stateTransition = 11'd463;
      4: stateTransition = 11'd463;
      5: stateTransition = 11'd463;
      6: stateTransition = 11'd463;
      7: stateTransition = 11'd463;
      8: stateTransition = 11'd463;
      9: stateTransition = 11'd463;
      10: stateTransition = 11'd463;
      11: stateTransition = 11'd463;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd463;
      14: stateTransition = 11'd463;
      15: stateTransition = 11'd463;
      16: stateTransition = 11'd463;
      default: stateTransition = 11'bX;
    endcase
    464: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd464;
      2: stateTransition = 11'd464;
      3: stateTransition = 11'd464;
      4: stateTransition = 11'd464;
      5: stateTransition = 11'd464;
      6: stateTransition = 11'd464;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd464;
      9: stateTransition = 11'd464;
      10: stateTransition = 11'd464;
      11: stateTransition = 11'd464;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd464;
      14: stateTransition = 11'd464;
      15: stateTransition = 11'd464;
      16: stateTransition = 11'd464;
      default: stateTransition = 11'bX;
    endcase
    465: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd465;
      2: stateTransition = 11'd465;
      3: stateTransition = 11'd465;
      4: stateTransition = 11'd465;
      5: stateTransition = 11'd465;
      6: stateTransition = 11'd465;
      7: stateTransition = 11'd465;
      8: stateTransition = 11'd465;
      9: stateTransition = 11'd465;
      10: stateTransition = 11'd465;
      11: stateTransition = 11'd465;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd465;
      14: stateTransition = 11'd465;
      15: stateTransition = 11'd465;
      16: stateTransition = 11'd465;
      default: stateTransition = 11'bX;
    endcase
    466: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd466;
      5: stateTransition = 11'd466;
      6: stateTransition = 11'd466;
      7: stateTransition = 11'd466;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd466;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    467: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd467;
      2: stateTransition = 11'd467;
      3: stateTransition = 11'd467;
      4: stateTransition = 11'd467;
      5: stateTransition = 11'd467;
      6: stateTransition = 11'd467;
      7: stateTransition = 11'd467;
      8: stateTransition = 11'd467;
      9: stateTransition = 11'd467;
      10: stateTransition = 11'd467;
      11: stateTransition = 11'd467;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd467;
      14: stateTransition = 11'd467;
      15: stateTransition = 11'd467;
      16: stateTransition = 11'd467;
      default: stateTransition = 11'bX;
    endcase
    468: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd468;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd468;
      10: stateTransition = 11'd468;
      11: stateTransition = 11'd468;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd468;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd468;
      16: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    469: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd469;
      2: stateTransition = 11'd469;
      3: stateTransition = 11'd469;
      4: stateTransition = 11'd469;
      5: stateTransition = 11'd469;
      6: stateTransition = 11'd469;
      7: stateTransition = 11'd469;
      8: stateTransition = 11'd469;
      9: stateTransition = 11'd469;
      10: stateTransition = 11'd469;
      11: stateTransition = 11'd469;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd469;
      14: stateTransition = 11'd469;
      15: stateTransition = 11'd469;
      16: stateTransition = 11'd469;
      default: stateTransition = 11'bX;
    endcase
    470: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd470;
      2: stateTransition = 11'd470;
      3: stateTransition = 11'd470;
      4: stateTransition = 11'd470;
      5: stateTransition = 11'd470;
      6: stateTransition = 11'd470;
      7: stateTransition = 11'd470;
      8: stateTransition = 11'd470;
      9: stateTransition = 11'd470;
      10: stateTransition = 11'd470;
      11: stateTransition = 11'd470;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd470;
      14: stateTransition = 11'd470;
      15: stateTransition = 11'd470;
      16: stateTransition = 11'd470;
      default: stateTransition = 11'bX;
    endcase
    471: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd471;
      2: stateTransition = 11'd471;
      3: stateTransition = 11'd471;
      4: stateTransition = 11'd471;
      5: stateTransition = 11'd471;
      6: stateTransition = 11'd471;
      7: stateTransition = 11'd471;
      8: stateTransition = 11'd471;
      9: stateTransition = 11'd471;
      10: stateTransition = 11'd471;
      11: stateTransition = 11'd471;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd471;
      14: stateTransition = 11'd471;
      15: stateTransition = 11'd471;
      16: stateTransition = 11'd471;
      default: stateTransition = 11'bX;
    endcase
    472: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd472;
      2: stateTransition = 11'd472;
      3: stateTransition = 11'd472;
      4: stateTransition = 11'd472;
      5: stateTransition = 11'd472;
      6: stateTransition = 11'd472;
      7: stateTransition = 11'd472;
      8: stateTransition = 11'd472;
      9: stateTransition = 11'd472;
      10: stateTransition = 11'd472;
      11: stateTransition = 11'd472;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd472;
      14: stateTransition = 11'd472;
      15: stateTransition = 11'd472;
      16: stateTransition = 11'd472;
      default: stateTransition = 11'bX;
    endcase
    473: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd473;
      2: stateTransition = 11'd473;
      3: stateTransition = 11'd473;
      4: stateTransition = 11'd473;
      5: stateTransition = 11'd473;
      6: stateTransition = 11'd473;
      7: stateTransition = 11'd473;
      8: stateTransition = 11'd473;
      9: stateTransition = 11'd473;
      10: stateTransition = 11'd473;
      11: stateTransition = 11'd473;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd473;
      14: stateTransition = 11'd473;
      15: stateTransition = 11'd473;
      16: stateTransition = 11'd473;
      default: stateTransition = 11'bX;
    endcase
    474: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd474;
      2: stateTransition = 11'd474;
      3: stateTransition = 11'd474;
      4: stateTransition = 11'd474;
      5: stateTransition = 11'd474;
      6: stateTransition = 11'd474;
      7: stateTransition = 11'd474;
      8: stateTransition = 11'd474;
      9: stateTransition = 11'd474;
      10: stateTransition = 11'd474;
      11: stateTransition = 11'd474;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd474;
      14: stateTransition = 11'd474;
      15: stateTransition = 11'd474;
      16: stateTransition = 11'd474;
      default: stateTransition = 11'bX;
    endcase
    475: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd475;
      2: stateTransition = 11'd475;
      3: stateTransition = 11'd475;
      4: stateTransition = 11'd475;
      5: stateTransition = 11'd475;
      6: stateTransition = 11'd475;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd475;
      9: stateTransition = 11'd475;
      10: stateTransition = 11'd475;
      11: stateTransition = 11'd475;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd475;
      14: stateTransition = 11'd475;
      15: stateTransition = 11'd475;
      16: stateTransition = 11'd475;
      default: stateTransition = 11'bX;
    endcase
    476: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd476;
      5: stateTransition = 11'd476;
      6: stateTransition = 11'd476;
      7: stateTransition = 11'd476;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd476;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    477: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd477;
      2: stateTransition = 11'd477;
      3: stateTransition = 11'd477;
      4: stateTransition = 11'd477;
      5: stateTransition = 11'd477;
      6: stateTransition = 11'd477;
      7: stateTransition = 11'd477;
      8: stateTransition = 11'd477;
      9: stateTransition = 11'd477;
      10: stateTransition = 11'd477;
      11: stateTransition = 11'd477;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd477;
      14: stateTransition = 11'd477;
      15: stateTransition = 11'd477;
      16: stateTransition = 11'd477;
      default: stateTransition = 11'bX;
    endcase
    478: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd478;
      2: stateTransition = 11'd478;
      3: stateTransition = 11'd478;
      4: stateTransition = 11'd478;
      5: stateTransition = 11'd478;
      6: stateTransition = 11'd478;
      7: stateTransition = 11'd478;
      8: stateTransition = 11'd478;
      9: stateTransition = 11'd478;
      10: stateTransition = 11'd478;
      11: stateTransition = 11'd478;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd478;
      14: stateTransition = 11'd478;
      15: stateTransition = 11'd478;
      16: stateTransition = 11'd478;
      default: stateTransition = 11'bX;
    endcase
    479: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd479;
      2: stateTransition = 11'd479;
      3: stateTransition = 11'd479;
      4: stateTransition = 11'd479;
      5: stateTransition = 11'd479;
      6: stateTransition = 11'd479;
      7: stateTransition = 11'd479;
      8: stateTransition = 11'd479;
      9: stateTransition = 11'd479;
      10: stateTransition = 11'd479;
      11: stateTransition = 11'd479;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd479;
      14: stateTransition = 11'd479;
      15: stateTransition = 11'd479;
      16: stateTransition = 11'd479;
      default: stateTransition = 11'bX;
    endcase
    480: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd480;
      2: stateTransition = 11'd480;
      3: stateTransition = 11'd480;
      4: stateTransition = 11'd480;
      5: stateTransition = 11'd480;
      6: stateTransition = 11'd480;
      7: stateTransition = 11'd480;
      8: stateTransition = 11'd480;
      9: stateTransition = 11'd480;
      10: stateTransition = 11'd480;
      11: stateTransition = 11'd480;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd480;
      14: stateTransition = 11'd480;
      15: stateTransition = 11'd480;
      16: stateTransition = 11'd480;
      default: stateTransition = 11'bX;
    endcase
    481: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd481;
      2: stateTransition = 11'd481;
      3: stateTransition = 11'd481;
      4: stateTransition = 11'd481;
      5: stateTransition = 11'd481;
      6: stateTransition = 11'd481;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd481;
      9: stateTransition = 11'd481;
      10: stateTransition = 11'd481;
      11: stateTransition = 11'd481;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd481;
      14: stateTransition = 11'd481;
      15: stateTransition = 11'd481;
      16: stateTransition = 11'd481;
      default: stateTransition = 11'bX;
    endcase
    482: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd482;
      5: stateTransition = 11'd482;
      6: stateTransition = 11'd482;
      7: stateTransition = 11'd482;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd482;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    483: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd483;
      2: stateTransition = 11'd483;
      3: stateTransition = 11'd483;
      4: stateTransition = 11'd483;
      5: stateTransition = 11'd483;
      6: stateTransition = 11'd483;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd483;
      9: stateTransition = 11'd483;
      10: stateTransition = 11'd483;
      11: stateTransition = 11'd483;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd483;
      14: stateTransition = 11'd483;
      15: stateTransition = 11'd483;
      16: stateTransition = 11'd483;
      default: stateTransition = 11'bX;
    endcase
    484: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd484;
      2: stateTransition = 11'd484;
      3: stateTransition = 11'd484;
      4: stateTransition = 11'd484;
      5: stateTransition = 11'd484;
      6: stateTransition = 11'd484;
      7: stateTransition = 11'd484;
      8: stateTransition = 11'd484;
      9: stateTransition = 11'd484;
      10: stateTransition = 11'd484;
      11: stateTransition = 11'd484;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd484;
      14: stateTransition = 11'd484;
      15: stateTransition = 11'd484;
      16: stateTransition = 11'd484;
      default: stateTransition = 11'bX;
    endcase
    485: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd485;
      2: stateTransition = 11'd485;
      3: stateTransition = 11'd485;
      4: stateTransition = 11'd485;
      5: stateTransition = 11'd485;
      6: stateTransition = 11'd485;
      7: stateTransition = 11'd485;
      8: stateTransition = 11'd485;
      9: stateTransition = 11'd485;
      10: stateTransition = 11'd485;
      11: stateTransition = 11'd485;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd485;
      14: stateTransition = 11'd485;
      15: stateTransition = 11'd485;
      16: stateTransition = 11'd485;
      default: stateTransition = 11'bX;
    endcase
    486: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd486;
      2: stateTransition = 11'd486;
      3: stateTransition = 11'd486;
      4: stateTransition = 11'd486;
      5: stateTransition = 11'd486;
      6: stateTransition = 11'd486;
      7: stateTransition = 11'd486;
      8: stateTransition = 11'd486;
      9: stateTransition = 11'd486;
      10: stateTransition = 11'd486;
      11: stateTransition = 11'd486;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd486;
      14: stateTransition = 11'd486;
      15: stateTransition = 11'd486;
      16: stateTransition = 11'd486;
      default: stateTransition = 11'bX;
    endcase
    487: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd487;
      2: stateTransition = 11'd487;
      3: stateTransition = 11'd487;
      4: stateTransition = 11'd487;
      5: stateTransition = 11'd487;
      6: stateTransition = 11'd487;
      7: stateTransition = 11'd487;
      8: stateTransition = 11'd487;
      9: stateTransition = 11'd487;
      10: stateTransition = 11'd487;
      11: stateTransition = 11'd487;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd487;
      14: stateTransition = 11'd487;
      15: stateTransition = 11'd487;
      16: stateTransition = 11'd487;
      default: stateTransition = 11'bX;
    endcase
    488: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd488;
      2: stateTransition = 11'd488;
      3: stateTransition = 11'd488;
      4: stateTransition = 11'd488;
      5: stateTransition = 11'd488;
      6: stateTransition = 11'd488;
      7: stateTransition = 11'd488;
      8: stateTransition = 11'd488;
      9: stateTransition = 11'd488;
      10: stateTransition = 11'd488;
      11: stateTransition = 11'd488;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd488;
      14: stateTransition = 11'd488;
      15: stateTransition = 11'd488;
      16: stateTransition = 11'd488;
      default: stateTransition = 11'bX;
    endcase
    489: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd489;
      2: stateTransition = 11'd489;
      3: stateTransition = 11'd489;
      4: stateTransition = 11'd489;
      5: stateTransition = 11'd489;
      6: stateTransition = 11'd489;
      7: stateTransition = 11'd489;
      8: stateTransition = 11'd489;
      9: stateTransition = 11'd489;
      10: stateTransition = 11'd489;
      11: stateTransition = 11'd489;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd489;
      14: stateTransition = 11'd489;
      15: stateTransition = 11'd489;
      16: stateTransition = 11'd489;
      default: stateTransition = 11'bX;
    endcase
    490: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd490;
      2: stateTransition = 11'd490;
      3: stateTransition = 11'd490;
      4: stateTransition = 11'd490;
      5: stateTransition = 11'd490;
      6: stateTransition = 11'd490;
      7: stateTransition = 11'd490;
      8: stateTransition = 11'd490;
      9: stateTransition = 11'd490;
      10: stateTransition = 11'd490;
      11: stateTransition = 11'd490;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd490;
      14: stateTransition = 11'd490;
      15: stateTransition = 11'd490;
      16: stateTransition = 11'd490;
      default: stateTransition = 11'bX;
    endcase
    491: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd491;
      2: stateTransition = 11'd491;
      3: stateTransition = 11'd491;
      4: stateTransition = 11'd491;
      5: stateTransition = 11'd491;
      6: stateTransition = 11'd491;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd491;
      9: stateTransition = 11'd491;
      10: stateTransition = 11'd491;
      11: stateTransition = 11'd491;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd491;
      14: stateTransition = 11'd491;
      15: stateTransition = 11'd491;
      16: stateTransition = 11'd491;
      default: stateTransition = 11'bX;
    endcase
    492: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd492;
      2: stateTransition = 11'd492;
      3: stateTransition = 11'd492;
      4: stateTransition = 11'd492;
      5: stateTransition = 11'd492;
      6: stateTransition = 11'd492;
      7: stateTransition = 11'd492;
      8: stateTransition = 11'd492;
      9: stateTransition = 11'd492;
      10: stateTransition = 11'd492;
      11: stateTransition = 11'd492;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd492;
      14: stateTransition = 11'd492;
      15: stateTransition = 11'd492;
      16: stateTransition = 11'd492;
      default: stateTransition = 11'bX;
    endcase
    493: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd493;
      5: stateTransition = 11'd493;
      6: stateTransition = 11'd493;
      7: stateTransition = 11'd493;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd493;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    494: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd494;
      2: stateTransition = 11'd494;
      3: stateTransition = 11'd494;
      4: stateTransition = 11'd494;
      5: stateTransition = 11'd494;
      6: stateTransition = 11'd494;
      7: stateTransition = 11'd494;
      8: stateTransition = 11'd494;
      9: stateTransition = 11'd494;
      10: stateTransition = 11'd494;
      11: stateTransition = 11'd494;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd494;
      14: stateTransition = 11'd494;
      15: stateTransition = 11'd494;
      16: stateTransition = 11'd494;
      default: stateTransition = 11'bX;
    endcase
    495: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd495;
      2: stateTransition = 11'd495;
      3: stateTransition = 11'd495;
      4: stateTransition = 11'd495;
      5: stateTransition = 11'd495;
      6: stateTransition = 11'd495;
      7: stateTransition = 11'd495;
      8: stateTransition = 11'd495;
      9: stateTransition = 11'd495;
      10: stateTransition = 11'd495;
      11: stateTransition = 11'd495;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd495;
      14: stateTransition = 11'd495;
      15: stateTransition = 11'd495;
      16: stateTransition = 11'd495;
      default: stateTransition = 11'bX;
    endcase
    496: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd496;
      2: stateTransition = 11'd496;
      3: stateTransition = 11'd496;
      4: stateTransition = 11'd496;
      5: stateTransition = 11'd496;
      6: stateTransition = 11'd496;
      7: stateTransition = 11'd496;
      8: stateTransition = 11'd496;
      9: stateTransition = 11'd496;
      10: stateTransition = 11'd496;
      11: stateTransition = 11'd496;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd496;
      14: stateTransition = 11'd496;
      15: stateTransition = 11'd496;
      16: stateTransition = 11'd496;
      default: stateTransition = 11'bX;
    endcase
    497: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd497;
      2: stateTransition = 11'd497;
      3: stateTransition = 11'd497;
      4: stateTransition = 11'd497;
      5: stateTransition = 11'd497;
      6: stateTransition = 11'd497;
      7: stateTransition = 11'd497;
      8: stateTransition = 11'd497;
      9: stateTransition = 11'd497;
      10: stateTransition = 11'd497;
      11: stateTransition = 11'd497;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd497;
      14: stateTransition = 11'd497;
      15: stateTransition = 11'd497;
      16: stateTransition = 11'd497;
      default: stateTransition = 11'bX;
    endcase
    498: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd498;
      2: stateTransition = 11'd498;
      3: stateTransition = 11'd498;
      4: stateTransition = 11'd498;
      5: stateTransition = 11'd498;
      6: stateTransition = 11'd498;
      7: stateTransition = 11'd498;
      8: stateTransition = 11'd498;
      9: stateTransition = 11'd498;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd498;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd498;
      14: stateTransition = 11'd498;
      15: stateTransition = 11'd498;
      16: stateTransition = 11'd498;
      default: stateTransition = 11'bX;
    endcase
    499: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd499;
      2: stateTransition = 11'd499;
      3: stateTransition = 11'd499;
      4: stateTransition = 11'd499;
      5: stateTransition = 11'd499;
      6: stateTransition = 11'd499;
      7: stateTransition = 11'd499;
      8: stateTransition = 11'd499;
      9: stateTransition = 11'd499;
      10: stateTransition = 11'd499;
      11: stateTransition = 11'd499;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd499;
      14: stateTransition = 11'd499;
      15: stateTransition = 11'd499;
      16: stateTransition = 11'd499;
      default: stateTransition = 11'bX;
    endcase
    500: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd500;
      5: stateTransition = 11'd500;
      6: stateTransition = 11'd500;
      7: stateTransition = 11'd500;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd500;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    501: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd501;
      2: stateTransition = 11'd501;
      3: stateTransition = 11'd501;
      4: stateTransition = 11'd501;
      5: stateTransition = 11'd501;
      6: stateTransition = 11'd501;
      7: stateTransition = 11'd501;
      8: stateTransition = 11'd501;
      9: stateTransition = 11'd501;
      10: stateTransition = 11'd501;
      11: stateTransition = 11'd501;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd501;
      14: stateTransition = 11'd501;
      15: stateTransition = 11'd501;
      16: stateTransition = 11'd501;
      default: stateTransition = 11'bX;
    endcase
    502: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd502;
      2: stateTransition = 11'd502;
      3: stateTransition = 11'd502;
      4: stateTransition = 11'd502;
      5: stateTransition = 11'd502;
      6: stateTransition = 11'd502;
      7: stateTransition = 11'd502;
      8: stateTransition = 11'd502;
      9: stateTransition = 11'd502;
      10: stateTransition = 11'd502;
      11: stateTransition = 11'd502;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd502;
      14: stateTransition = 11'd502;
      15: stateTransition = 11'd502;
      16: stateTransition = 11'd502;
      default: stateTransition = 11'bX;
    endcase
    503: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd503;
      5: stateTransition = 11'd503;
      6: stateTransition = 11'd503;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd503;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    504: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd504;
      2: stateTransition = 11'd504;
      3: stateTransition = 11'd504;
      4: stateTransition = 11'd504;
      5: stateTransition = 11'd504;
      6: stateTransition = 11'd504;
      7: stateTransition = 11'd504;
      8: stateTransition = 11'd504;
      9: stateTransition = 11'd504;
      10: stateTransition = 11'd504;
      11: stateTransition = 11'd504;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd504;
      14: stateTransition = 11'd504;
      15: stateTransition = 11'd504;
      16: stateTransition = 11'd504;
      default: stateTransition = 11'bX;
    endcase
    505: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd505;
      2: stateTransition = 11'd505;
      3: stateTransition = 11'd505;
      4: stateTransition = 11'd505;
      5: stateTransition = 11'd505;
      6: stateTransition = 11'd505;
      7: stateTransition = 11'd505;
      8: stateTransition = 11'd505;
      9: stateTransition = 11'd505;
      10: stateTransition = 11'd505;
      11: stateTransition = 11'd505;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd505;
      14: stateTransition = 11'd505;
      15: stateTransition = 11'd505;
      16: stateTransition = 11'd505;
      default: stateTransition = 11'bX;
    endcase
    506: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd506;
      2: stateTransition = 11'd506;
      3: stateTransition = 11'd506;
      4: stateTransition = 11'd506;
      5: stateTransition = 11'd506;
      6: stateTransition = 11'd506;
      7: stateTransition = 11'd506;
      8: stateTransition = 11'd506;
      9: stateTransition = 11'd506;
      10: stateTransition = 11'd506;
      11: stateTransition = 11'd506;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd506;
      14: stateTransition = 11'd506;
      15: stateTransition = 11'd506;
      16: stateTransition = 11'd506;
      default: stateTransition = 11'bX;
    endcase
    507: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd507;
      2: stateTransition = 11'd507;
      3: stateTransition = 11'd507;
      4: stateTransition = 11'd507;
      5: stateTransition = 11'd507;
      6: stateTransition = 11'd507;
      7: stateTransition = 11'd507;
      8: stateTransition = 11'd507;
      9: stateTransition = 11'd507;
      10: stateTransition = 11'd507;
      11: stateTransition = 11'd507;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd507;
      14: stateTransition = 11'd507;
      15: stateTransition = 11'd507;
      16: stateTransition = 11'd507;
      default: stateTransition = 11'bX;
    endcase
    508: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd508;
      2: stateTransition = 11'd508;
      3: stateTransition = 11'd508;
      4: stateTransition = 11'd508;
      5: stateTransition = 11'd508;
      6: stateTransition = 11'd508;
      7: stateTransition = 11'd508;
      8: stateTransition = 11'd508;
      9: stateTransition = 11'd508;
      10: stateTransition = 11'd508;
      11: stateTransition = 11'd508;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd508;
      14: stateTransition = 11'd508;
      15: stateTransition = 11'd508;
      16: stateTransition = 11'd508;
      default: stateTransition = 11'bX;
    endcase
    509: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd509;
      2: stateTransition = 11'd509;
      3: stateTransition = 11'd509;
      4: stateTransition = 11'd509;
      5: stateTransition = 11'd509;
      6: stateTransition = 11'd509;
      7: stateTransition = 11'd509;
      8: stateTransition = 11'd509;
      9: stateTransition = 11'd509;
      10: stateTransition = 11'd509;
      11: stateTransition = 11'd509;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd509;
      14: stateTransition = 11'd509;
      15: stateTransition = 11'd509;
      16: stateTransition = 11'd509;
      default: stateTransition = 11'bX;
    endcase
    510: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd510;
      2: stateTransition = 11'd510;
      3: stateTransition = 11'd510;
      4: stateTransition = 11'd510;
      5: stateTransition = 11'd510;
      6: stateTransition = 11'd510;
      7: stateTransition = 11'd510;
      8: stateTransition = 11'd510;
      9: stateTransition = 11'd510;
      10: stateTransition = 11'd510;
      11: stateTransition = 11'd510;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd510;
      14: stateTransition = 11'd510;
      15: stateTransition = 11'd510;
      16: stateTransition = 11'd510;
      default: stateTransition = 11'bX;
    endcase
    511: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd511;
      2: stateTransition = 11'd511;
      3: stateTransition = 11'd511;
      4: stateTransition = 11'd511;
      5: stateTransition = 11'd511;
      6: stateTransition = 11'd511;
      7: stateTransition = 11'd511;
      8: stateTransition = 11'd511;
      9: stateTransition = 11'd511;
      10: stateTransition = 11'd511;
      11: stateTransition = 11'd511;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd511;
      14: stateTransition = 11'd511;
      15: stateTransition = 11'd511;
      16: stateTransition = 11'd511;
      default: stateTransition = 11'bX;
    endcase
    512: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd512;
      2: stateTransition = 11'd512;
      3: stateTransition = 11'd512;
      4: stateTransition = 11'd512;
      5: stateTransition = 11'd512;
      6: stateTransition = 11'd512;
      7: stateTransition = 11'd512;
      8: stateTransition = 11'd512;
      9: stateTransition = 11'd512;
      10: stateTransition = 11'd512;
      11: stateTransition = 11'd512;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd512;
      14: stateTransition = 11'd512;
      15: stateTransition = 11'd512;
      16: stateTransition = 11'd512;
      default: stateTransition = 11'bX;
    endcase
    513: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd513;
      2: stateTransition = 11'd513;
      3: stateTransition = 11'd513;
      4: stateTransition = 11'd513;
      5: stateTransition = 11'd513;
      6: stateTransition = 11'd513;
      7: stateTransition = 11'd513;
      8: stateTransition = 11'd513;
      9: stateTransition = 11'd513;
      10: stateTransition = 11'd513;
      11: stateTransition = 11'd513;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd513;
      14: stateTransition = 11'd513;
      15: stateTransition = 11'd513;
      16: stateTransition = 11'd513;
      default: stateTransition = 11'bX;
    endcase
    514: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd514;
      2: stateTransition = 11'd514;
      3: stateTransition = 11'd514;
      4: stateTransition = 11'd514;
      5: stateTransition = 11'd514;
      6: stateTransition = 11'd514;
      7: stateTransition = 11'd514;
      8: stateTransition = 11'd514;
      9: stateTransition = 11'd514;
      10: stateTransition = 11'd514;
      11: stateTransition = 11'd514;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd514;
      14: stateTransition = 11'd514;
      15: stateTransition = 11'd514;
      16: stateTransition = 11'd514;
      default: stateTransition = 11'bX;
    endcase
    515: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd515;
      2: stateTransition = 11'd515;
      3: stateTransition = 11'd515;
      4: stateTransition = 11'd515;
      5: stateTransition = 11'd515;
      6: stateTransition = 11'd515;
      7: stateTransition = 11'd515;
      8: stateTransition = 11'd515;
      9: stateTransition = 11'd515;
      10: stateTransition = 11'd515;
      11: stateTransition = 11'd515;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd515;
      14: stateTransition = 11'd515;
      15: stateTransition = 11'd515;
      16: stateTransition = 11'd515;
      default: stateTransition = 11'bX;
    endcase
    516: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd516;
      2: stateTransition = 11'd516;
      3: stateTransition = 11'd516;
      4: stateTransition = 11'd516;
      5: stateTransition = 11'd516;
      6: stateTransition = 11'd516;
      7: stateTransition = 11'd516;
      8: stateTransition = 11'd516;
      9: stateTransition = 11'd516;
      10: stateTransition = 11'd516;
      11: stateTransition = 11'd516;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd516;
      14: stateTransition = 11'd516;
      15: stateTransition = 11'd516;
      16: stateTransition = 11'd516;
      default: stateTransition = 11'bX;
    endcase
    517: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd517;
      2: stateTransition = 11'd517;
      3: stateTransition = 11'd517;
      4: stateTransition = 11'd517;
      5: stateTransition = 11'd517;
      6: stateTransition = 11'd517;
      7: stateTransition = 11'd517;
      8: stateTransition = 11'd517;
      9: stateTransition = 11'd517;
      10: stateTransition = 11'd517;
      11: stateTransition = 11'd517;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd517;
      14: stateTransition = 11'd517;
      15: stateTransition = 11'd517;
      16: stateTransition = 11'd517;
      default: stateTransition = 11'bX;
    endcase
    518: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd518;
      2: stateTransition = 11'd518;
      3: stateTransition = 11'd518;
      4: stateTransition = 11'd518;
      5: stateTransition = 11'd518;
      6: stateTransition = 11'd518;
      7: stateTransition = 11'd518;
      8: stateTransition = 11'd518;
      9: stateTransition = 11'd518;
      10: stateTransition = 11'd518;
      11: stateTransition = 11'd518;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd518;
      14: stateTransition = 11'd518;
      15: stateTransition = 11'd518;
      16: stateTransition = 11'd518;
      default: stateTransition = 11'bX;
    endcase
    519: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd519;
      2: stateTransition = 11'd519;
      3: stateTransition = 11'd519;
      4: stateTransition = 11'd519;
      5: stateTransition = 11'd519;
      6: stateTransition = 11'd519;
      7: stateTransition = 11'd519;
      8: stateTransition = 11'd519;
      9: stateTransition = 11'd519;
      10: stateTransition = 11'd519;
      11: stateTransition = 11'd519;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd519;
      14: stateTransition = 11'd519;
      15: stateTransition = 11'd519;
      16: stateTransition = 11'd519;
      default: stateTransition = 11'bX;
    endcase
    520: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd520;
      2: stateTransition = 11'd520;
      3: stateTransition = 11'd520;
      4: stateTransition = 11'd520;
      5: stateTransition = 11'd520;
      6: stateTransition = 11'd520;
      7: stateTransition = 11'd520;
      8: stateTransition = 11'd520;
      9: stateTransition = 11'd520;
      10: stateTransition = 11'd520;
      11: stateTransition = 11'd520;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd520;
      14: stateTransition = 11'd520;
      15: stateTransition = 11'd520;
      16: stateTransition = 11'd520;
      default: stateTransition = 11'bX;
    endcase
    521: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd521;
      2: stateTransition = 11'd521;
      3: stateTransition = 11'd521;
      4: stateTransition = 11'd521;
      5: stateTransition = 11'd521;
      6: stateTransition = 11'd521;
      7: stateTransition = 11'd521;
      8: stateTransition = 11'd521;
      9: stateTransition = 11'd521;
      10: stateTransition = 11'd521;
      11: stateTransition = 11'd521;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd521;
      14: stateTransition = 11'd521;
      15: stateTransition = 11'd521;
      16: stateTransition = 11'd521;
      default: stateTransition = 11'bX;
    endcase
    522: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd522;
      2: stateTransition = 11'd522;
      3: stateTransition = 11'd522;
      4: stateTransition = 11'd522;
      5: stateTransition = 11'd522;
      6: stateTransition = 11'd522;
      7: stateTransition = 11'd522;
      8: stateTransition = 11'd522;
      9: stateTransition = 11'd522;
      10: stateTransition = 11'd522;
      11: stateTransition = 11'd522;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd522;
      14: stateTransition = 11'd522;
      15: stateTransition = 11'd522;
      16: stateTransition = 11'd522;
      default: stateTransition = 11'bX;
    endcase
    523: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd523;
      2: stateTransition = 11'd523;
      3: stateTransition = 11'd523;
      4: stateTransition = 11'd523;
      5: stateTransition = 11'd523;
      6: stateTransition = 11'd523;
      7: stateTransition = 11'd523;
      8: stateTransition = 11'd523;
      9: stateTransition = 11'd523;
      10: stateTransition = 11'd523;
      11: stateTransition = 11'd523;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd523;
      14: stateTransition = 11'd523;
      15: stateTransition = 11'd523;
      16: stateTransition = 11'd523;
      default: stateTransition = 11'bX;
    endcase
    524: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd524;
      2: stateTransition = 11'd524;
      3: stateTransition = 11'd524;
      4: stateTransition = 11'd524;
      5: stateTransition = 11'd524;
      6: stateTransition = 11'd524;
      7: stateTransition = 11'd524;
      8: stateTransition = 11'd524;
      9: stateTransition = 11'd524;
      10: stateTransition = 11'd524;
      11: stateTransition = 11'd524;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd524;
      14: stateTransition = 11'd524;
      15: stateTransition = 11'd524;
      16: stateTransition = 11'd524;
      default: stateTransition = 11'bX;
    endcase
    525: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd525;
      2: stateTransition = 11'd525;
      3: stateTransition = 11'd525;
      4: stateTransition = 11'd525;
      5: stateTransition = 11'd525;
      6: stateTransition = 11'd525;
      7: stateTransition = 11'd525;
      8: stateTransition = 11'd525;
      9: stateTransition = 11'd525;
      10: stateTransition = 11'd525;
      11: stateTransition = 11'd525;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd525;
      14: stateTransition = 11'd525;
      15: stateTransition = 11'd525;
      16: stateTransition = 11'd525;
      default: stateTransition = 11'bX;
    endcase
    526: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd526;
      2: stateTransition = 11'd526;
      3: stateTransition = 11'd526;
      4: stateTransition = 11'd526;
      5: stateTransition = 11'd526;
      6: stateTransition = 11'd526;
      7: stateTransition = 11'd526;
      8: stateTransition = 11'd526;
      9: stateTransition = 11'd526;
      10: stateTransition = 11'd526;
      11: stateTransition = 11'd526;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd526;
      14: stateTransition = 11'd526;
      15: stateTransition = 11'd526;
      16: stateTransition = 11'd526;
      default: stateTransition = 11'bX;
    endcase
    527: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd527;
      2: stateTransition = 11'd527;
      3: stateTransition = 11'd527;
      4: stateTransition = 11'd527;
      5: stateTransition = 11'd527;
      6: stateTransition = 11'd527;
      7: stateTransition = 11'd527;
      8: stateTransition = 11'd527;
      9: stateTransition = 11'd527;
      10: stateTransition = 11'd527;
      11: stateTransition = 11'd527;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd527;
      14: stateTransition = 11'd527;
      15: stateTransition = 11'd527;
      16: stateTransition = 11'd527;
      default: stateTransition = 11'bX;
    endcase
    528: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd528;
      2: stateTransition = 11'd528;
      3: stateTransition = 11'd528;
      4: stateTransition = 11'd528;
      5: stateTransition = 11'd528;
      6: stateTransition = 11'd528;
      7: stateTransition = 11'd528;
      8: stateTransition = 11'd528;
      9: stateTransition = 11'd528;
      10: stateTransition = 11'd528;
      11: stateTransition = 11'd528;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd528;
      14: stateTransition = 11'd528;
      15: stateTransition = 11'd528;
      16: stateTransition = 11'd528;
      default: stateTransition = 11'bX;
    endcase
    529: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd529;
      2: stateTransition = 11'd529;
      3: stateTransition = 11'd529;
      4: stateTransition = 11'd529;
      5: stateTransition = 11'd529;
      6: stateTransition = 11'd529;
      7: stateTransition = 11'd529;
      8: stateTransition = 11'd529;
      9: stateTransition = 11'd529;
      10: stateTransition = 11'd529;
      11: stateTransition = 11'd529;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd529;
      14: stateTransition = 11'd529;
      15: stateTransition = 11'd529;
      16: stateTransition = 11'd529;
      default: stateTransition = 11'bX;
    endcase
    530: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd530;
      2: stateTransition = 11'd530;
      3: stateTransition = 11'd530;
      4: stateTransition = 11'd530;
      5: stateTransition = 11'd530;
      6: stateTransition = 11'd530;
      7: stateTransition = 11'd530;
      8: stateTransition = 11'd530;
      9: stateTransition = 11'd530;
      10: stateTransition = 11'd530;
      11: stateTransition = 11'd530;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd530;
      14: stateTransition = 11'd530;
      15: stateTransition = 11'd530;
      16: stateTransition = 11'd530;
      default: stateTransition = 11'bX;
    endcase
    531: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd531;
      2: stateTransition = 11'd531;
      3: stateTransition = 11'd531;
      4: stateTransition = 11'd531;
      5: stateTransition = 11'd531;
      6: stateTransition = 11'd531;
      7: stateTransition = 11'd531;
      8: stateTransition = 11'd531;
      9: stateTransition = 11'd531;
      10: stateTransition = 11'd531;
      11: stateTransition = 11'd531;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd531;
      14: stateTransition = 11'd531;
      15: stateTransition = 11'd531;
      16: stateTransition = 11'd531;
      default: stateTransition = 11'bX;
    endcase
    532: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd532;
      2: stateTransition = 11'd532;
      3: stateTransition = 11'd532;
      4: stateTransition = 11'd532;
      5: stateTransition = 11'd532;
      6: stateTransition = 11'd532;
      7: stateTransition = 11'd532;
      8: stateTransition = 11'd532;
      9: stateTransition = 11'd532;
      10: stateTransition = 11'd532;
      11: stateTransition = 11'd532;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd532;
      14: stateTransition = 11'd532;
      15: stateTransition = 11'd532;
      16: stateTransition = 11'd532;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
