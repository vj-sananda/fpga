`timescale 1ns/1ps

`define ENABLED_REGEX_CATEGORY_dns TRUE

module CATEGORY_dns_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_CATEGORY_dns

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd1;
    1: charMap = 8'd2;
    2: charMap = 8'd7;
    3: charMap = 8'd35;
    4: charMap = 8'd35;
    5: charMap = 8'd8;
    6: charMap = 8'd8;
    7: charMap = 8'd34;
    8: charMap = 8'd34;
    9: charMap = 8'd34;
    10: charMap = 8'd4;
    11: charMap = 8'd34;
    12: charMap = 8'd34;
    13: charMap = 8'd4;
    14: charMap = 8'd34;
    15: charMap = 8'd34;
    16: charMap = 8'd34;
    17: charMap = 8'd3;
    18: charMap = 8'd3;
    19: charMap = 8'd3;
    20: charMap = 8'd3;
    21: charMap = 8'd3;
    22: charMap = 8'd3;
    23: charMap = 8'd3;
    24: charMap = 8'd3;
    25: charMap = 8'd3;
    26: charMap = 8'd3;
    27: charMap = 8'd3;
    28: charMap = 8'd3;
    29: charMap = 8'd3;
    30: charMap = 8'd3;
    31: charMap = 8'd3;
    32: charMap = 8'd3;
    33: charMap = 8'd3;
    34: charMap = 8'd3;
    35: charMap = 8'd3;
    36: charMap = 8'd3;
    37: charMap = 8'd3;
    38: charMap = 8'd3;
    39: charMap = 8'd3;
    40: charMap = 8'd3;
    41: charMap = 8'd3;
    42: charMap = 8'd3;
    43: charMap = 8'd3;
    44: charMap = 8'd3;
    45: charMap = 8'd3;
    46: charMap = 8'd3;
    47: charMap = 8'd3;
    48: charMap = 8'd5;
    49: charMap = 8'd5;
    50: charMap = 8'd5;
    51: charMap = 8'd5;
    52: charMap = 8'd5;
    53: charMap = 8'd5;
    54: charMap = 8'd5;
    55: charMap = 8'd5;
    56: charMap = 8'd5;
    57: charMap = 8'd5;
    58: charMap = 8'd3;
    59: charMap = 8'd3;
    60: charMap = 8'd3;
    61: charMap = 8'd3;
    62: charMap = 8'd3;
    63: charMap = 8'd3;
    64: charMap = 8'd1;
    65: charMap = 8'd1;
    66: charMap = 8'd1;
    67: charMap = 8'd1;
    68: charMap = 8'd1;
    69: charMap = 8'd1;
    70: charMap = 8'd1;
    71: charMap = 8'd1;
    72: charMap = 8'd1;
    73: charMap = 8'd1;
    74: charMap = 8'd1;
    75: charMap = 8'd1;
    76: charMap = 8'd1;
    77: charMap = 8'd1;
    78: charMap = 8'd1;
    79: charMap = 8'd1;
    80: charMap = 8'd1;
    81: charMap = 8'd1;
    82: charMap = 8'd1;
    83: charMap = 8'd1;
    84: charMap = 8'd1;
    85: charMap = 8'd1;
    86: charMap = 8'd1;
    87: charMap = 8'd1;
    88: charMap = 8'd1;
    89: charMap = 8'd1;
    90: charMap = 8'd1;
    91: charMap = 8'd1;
    92: charMap = 8'd1;
    93: charMap = 8'd1;
    94: charMap = 8'd1;
    95: charMap = 8'd1;
    96: charMap = 8'd1;
    97: charMap = 8'd9;
    98: charMap = 8'd14;
    99: charMap = 8'd17;
    100: charMap = 8'd19;
    101: charMap = 8'd10;
    102: charMap = 8'd24;
    103: charMap = 8'd21;
    104: charMap = 8'd30;
    105: charMap = 8'd15;
    106: charMap = 8'd31;
    107: charMap = 8'd33;
    108: charMap = 8'd26;
    109: charMap = 8'd18;
    110: charMap = 8'd23;
    111: charMap = 8'd12;
    112: charMap = 8'd13;
    113: charMap = 8'd28;
    114: charMap = 8'd11;
    115: charMap = 8'd27;
    116: charMap = 8'd25;
    117: charMap = 8'd20;
    118: charMap = 8'd22;
    119: charMap = 8'd29;
    120: charMap = 8'd6;
    121: charMap = 8'd32;
    122: charMap = 8'd16;
    123: charMap = 8'd1;
    124: charMap = 8'd1;
    125: charMap = 8'd1;
    126: charMap = 8'd1;
    127: charMap = 8'd1;
    128: charMap = 8'd1;
    129: charMap = 8'd1;
    130: charMap = 8'd1;
    131: charMap = 8'd1;
    132: charMap = 8'd1;
    133: charMap = 8'd1;
    134: charMap = 8'd1;
    135: charMap = 8'd1;
    136: charMap = 8'd1;
    137: charMap = 8'd1;
    138: charMap = 8'd1;
    139: charMap = 8'd1;
    140: charMap = 8'd1;
    141: charMap = 8'd1;
    142: charMap = 8'd1;
    143: charMap = 8'd1;
    144: charMap = 8'd1;
    145: charMap = 8'd1;
    146: charMap = 8'd1;
    147: charMap = 8'd1;
    148: charMap = 8'd1;
    149: charMap = 8'd1;
    150: charMap = 8'd1;
    151: charMap = 8'd1;
    152: charMap = 8'd1;
    153: charMap = 8'd1;
    154: charMap = 8'd1;
    155: charMap = 8'd1;
    156: charMap = 8'd1;
    157: charMap = 8'd1;
    158: charMap = 8'd1;
    159: charMap = 8'd1;
    160: charMap = 8'd1;
    161: charMap = 8'd1;
    162: charMap = 8'd1;
    163: charMap = 8'd1;
    164: charMap = 8'd1;
    165: charMap = 8'd1;
    166: charMap = 8'd1;
    167: charMap = 8'd1;
    168: charMap = 8'd1;
    169: charMap = 8'd1;
    170: charMap = 8'd1;
    171: charMap = 8'd1;
    172: charMap = 8'd1;
    173: charMap = 8'd1;
    174: charMap = 8'd1;
    175: charMap = 8'd1;
    176: charMap = 8'd1;
    177: charMap = 8'd1;
    178: charMap = 8'd1;
    179: charMap = 8'd1;
    180: charMap = 8'd1;
    181: charMap = 8'd1;
    182: charMap = 8'd1;
    183: charMap = 8'd1;
    184: charMap = 8'd1;
    185: charMap = 8'd1;
    186: charMap = 8'd1;
    187: charMap = 8'd1;
    188: charMap = 8'd1;
    189: charMap = 8'd1;
    190: charMap = 8'd1;
    191: charMap = 8'd1;
    192: charMap = 8'd1;
    193: charMap = 8'd1;
    194: charMap = 8'd1;
    195: charMap = 8'd1;
    196: charMap = 8'd1;
    197: charMap = 8'd1;
    198: charMap = 8'd1;
    199: charMap = 8'd1;
    200: charMap = 8'd1;
    201: charMap = 8'd1;
    202: charMap = 8'd1;
    203: charMap = 8'd1;
    204: charMap = 8'd1;
    205: charMap = 8'd1;
    206: charMap = 8'd1;
    207: charMap = 8'd1;
    208: charMap = 8'd1;
    209: charMap = 8'd1;
    210: charMap = 8'd1;
    211: charMap = 8'd1;
    212: charMap = 8'd1;
    213: charMap = 8'd1;
    214: charMap = 8'd1;
    215: charMap = 8'd1;
    216: charMap = 8'd1;
    217: charMap = 8'd1;
    218: charMap = 8'd1;
    219: charMap = 8'd1;
    220: charMap = 8'd1;
    221: charMap = 8'd1;
    222: charMap = 8'd1;
    223: charMap = 8'd1;
    224: charMap = 8'd1;
    225: charMap = 8'd1;
    226: charMap = 8'd1;
    227: charMap = 8'd1;
    228: charMap = 8'd1;
    229: charMap = 8'd1;
    230: charMap = 8'd1;
    231: charMap = 8'd1;
    232: charMap = 8'd1;
    233: charMap = 8'd1;
    234: charMap = 8'd1;
    235: charMap = 8'd1;
    236: charMap = 8'd1;
    237: charMap = 8'd1;
    238: charMap = 8'd1;
    239: charMap = 8'd1;
    240: charMap = 8'd1;
    241: charMap = 8'd1;
    242: charMap = 8'd1;
    243: charMap = 8'd1;
    244: charMap = 8'd1;
    245: charMap = 8'd1;
    246: charMap = 8'd1;
    247: charMap = 8'd1;
    248: charMap = 8'd1;
    249: charMap = 8'd1;
    250: charMap = 8'd1;
    251: charMap = 8'd1;
    252: charMap = 8'd1;
    253: charMap = 8'd1;
    254: charMap = 8'd1;
    255: charMap = 8'd36;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd2;
    3: stateMap = 11'd3;
    4: stateMap = 11'd4;
    5: stateMap = 11'd5;
    6: stateMap = 11'd1;
    7: stateMap = 11'd6;
    8: stateMap = 11'd7;
    9: stateMap = 11'd8;
    10: stateMap = 11'd9;
    11: stateMap = 11'd10;
    12: stateMap = 11'd11;
    13: stateMap = 11'd4;
    14: stateMap = 11'd12;
    15: stateMap = 11'd13;
    16: stateMap = 11'd14;
    17: stateMap = 11'd15;
    18: stateMap = 11'd16;
    19: stateMap = 11'd17;
    20: stateMap = 11'd18;
    21: stateMap = 11'd19;
    22: stateMap = 11'd20;
    23: stateMap = 11'd21;
    24: stateMap = 11'd22;
    25: stateMap = 11'd23;
    26: stateMap = 11'd24;
    27: stateMap = 11'd25;
    28: stateMap = 11'd26;
    29: stateMap = 11'd27;
    30: stateMap = 11'd7;
    31: stateMap = 11'd28;
    32: stateMap = 11'd29;
    33: stateMap = 11'd30;
    34: stateMap = 11'd31;
    35: stateMap = 11'd32;
    36: stateMap = 11'd33;
    37: stateMap = 11'd34;
    38: stateMap = 11'd35;
    39: stateMap = 11'd36;
    40: stateMap = 11'd37;
    41: stateMap = 11'd38;
    42: stateMap = 11'd39;
    43: stateMap = 11'd40;
    44: stateMap = 11'd41;
    45: stateMap = 11'd42;
    46: stateMap = 11'd43;
    47: stateMap = 11'd44;
    48: stateMap = 11'd45;
    49: stateMap = 11'd46;
    50: stateMap = 11'd47;
    51: stateMap = 11'd48;
    52: stateMap = 11'd49;
    53: stateMap = 11'd50;
    54: stateMap = 11'd51;
    55: stateMap = 11'd52;
    56: stateMap = 11'd53;
    57: stateMap = 11'd54;
    58: stateMap = 11'd55;
    59: stateMap = 11'd56;
    60: stateMap = 11'd57;
    61: stateMap = 11'd58;
    62: stateMap = 11'd59;
    63: stateMap = 11'd60;
    64: stateMap = 11'd54;
    65: stateMap = 11'd61;
    66: stateMap = 11'd62;
    67: stateMap = 11'd63;
    68: stateMap = 11'd64;
    69: stateMap = 11'd65;
    70: stateMap = 11'd66;
    71: stateMap = 11'd67;
    72: stateMap = 11'd68;
    73: stateMap = 11'd2;
    74: stateMap = 11'd69;
    75: stateMap = 11'd70;
    76: stateMap = 11'd71;
    77: stateMap = 11'd72;
    78: stateMap = 11'd73;
    79: stateMap = 11'd74;
    80: stateMap = 11'd75;
    81: stateMap = 11'd76;
    82: stateMap = 11'd77;
    83: stateMap = 11'd78;
    84: stateMap = 11'd79;
    85: stateMap = 11'd80;
    86: stateMap = 11'd81;
    87: stateMap = 11'd82;
    88: stateMap = 11'd83;
    89: stateMap = 11'd84;
    90: stateMap = 11'd85;
    91: stateMap = 11'd86;
    92: stateMap = 11'd87;
    93: stateMap = 11'd88;
    94: stateMap = 11'd89;
    95: stateMap = 11'd90;
    96: stateMap = 11'd91;
    97: stateMap = 11'd92;
    98: stateMap = 11'd93;
    99: stateMap = 11'd94;
    100: stateMap = 11'd95;
    101: stateMap = 11'd96;
    102: stateMap = 11'd97;
    103: stateMap = 11'd98;
    104: stateMap = 11'd99;
    105: stateMap = 11'd100;
    106: stateMap = 11'd101;
    107: stateMap = 11'd102;
    108: stateMap = 11'd103;
    109: stateMap = 11'd104;
    110: stateMap = 11'd105;
    111: stateMap = 11'd106;
    112: stateMap = 11'd107;
    113: stateMap = 11'd108;
    114: stateMap = 11'd109;
    115: stateMap = 11'd110;
    116: stateMap = 11'd111;
    117: stateMap = 11'd112;
    118: stateMap = 11'd113;
    119: stateMap = 11'd114;
    120: stateMap = 11'd115;
    121: stateMap = 11'd116;
    122: stateMap = 11'd117;
    123: stateMap = 11'd118;
    124: stateMap = 11'd119;
    125: stateMap = 11'd120;
    126: stateMap = 11'd121;
    127: stateMap = 11'd122;
    128: stateMap = 11'd123;
    129: stateMap = 11'd124;
    130: stateMap = 11'd125;
    131: stateMap = 11'd126;
    132: stateMap = 11'd127;
    133: stateMap = 11'd128;
    134: stateMap = 11'd129;
    135: stateMap = 11'd130;
    136: stateMap = 11'd131;
    137: stateMap = 11'd132;
    138: stateMap = 11'd133;
    139: stateMap = 11'd134;
    140: stateMap = 11'd135;
    141: stateMap = 11'd136;
    142: stateMap = 11'd41;
    143: stateMap = 11'd137;
    144: stateMap = 11'd138;
    145: stateMap = 11'd139;
    146: stateMap = 11'd140;
    147: stateMap = 11'd141;
    148: stateMap = 11'd142;
    149: stateMap = 11'd143;
    150: stateMap = 11'd144;
    151: stateMap = 11'd145;
    152: stateMap = 11'd146;
    153: stateMap = 11'd147;
    154: stateMap = 11'd148;
    155: stateMap = 11'd149;
    156: stateMap = 11'd150;
    157: stateMap = 11'd151;
    158: stateMap = 11'd152;
    159: stateMap = 11'd153;
    160: stateMap = 11'd154;
    161: stateMap = 11'd155;
    162: stateMap = 11'd156;
    163: stateMap = 11'd157;
    164: stateMap = 11'd158;
    165: stateMap = 11'd159;
    166: stateMap = 11'd160;
    167: stateMap = 11'd161;
    168: stateMap = 11'd162;
    169: stateMap = 11'd163;
    170: stateMap = 11'd164;
    171: stateMap = 11'd165;
    172: stateMap = 11'd166;
    173: stateMap = 11'd167;
    174: stateMap = 11'd168;
    175: stateMap = 11'd169;
    176: stateMap = 11'd170;
    177: stateMap = 11'd171;
    178: stateMap = 11'd172;
    179: stateMap = 11'd173;
    180: stateMap = 11'd174;
    181: stateMap = 11'd175;
    182: stateMap = 11'd176;
    183: stateMap = 11'd177;
    184: stateMap = 11'd178;
    185: stateMap = 11'd179;
    186: stateMap = 11'd180;
    187: stateMap = 11'd181;
    188: stateMap = 11'd182;
    189: stateMap = 11'd183;
    190: stateMap = 11'd184;
    191: stateMap = 11'd185;
    192: stateMap = 11'd186;
    193: stateMap = 11'd187;
    194: stateMap = 11'd188;
    195: stateMap = 11'd62;
    196: stateMap = 11'd189;
    197: stateMap = 11'd55;
    198: stateMap = 11'd59;
    199: stateMap = 11'd190;
    200: stateMap = 11'd191;
    201: stateMap = 11'd192;
    202: stateMap = 11'd193;
    203: stateMap = 11'd194;
    204: stateMap = 11'd195;
    205: stateMap = 11'd196;
    206: stateMap = 11'd197;
    207: stateMap = 11'd198;
    208: stateMap = 11'd199;
    209: stateMap = 11'd200;
    210: stateMap = 11'd201;
    211: stateMap = 11'd202;
    212: stateMap = 11'd203;
    213: stateMap = 11'd204;
    214: stateMap = 11'd205;
    215: stateMap = 11'd206;
    216: stateMap = 11'd207;
    217: stateMap = 11'd208;
    218: stateMap = 11'd209;
    219: stateMap = 11'd210;
    220: stateMap = 11'd211;
    221: stateMap = 11'd212;
    222: stateMap = 11'd213;
    223: stateMap = 11'd214;
    224: stateMap = 11'd215;
    225: stateMap = 11'd216;
    226: stateMap = 11'd217;
    227: stateMap = 11'd218;
    228: stateMap = 11'd219;
    229: stateMap = 11'd220;
    230: stateMap = 11'd221;
    231: stateMap = 11'd222;
    232: stateMap = 11'd223;
    233: stateMap = 11'd224;
    234: stateMap = 11'd225;
    235: stateMap = 11'd226;
    236: stateMap = 11'd227;
    237: stateMap = 11'd228;
    238: stateMap = 11'd229;
    239: stateMap = 11'd230;
    240: stateMap = 11'd231;
    241: stateMap = 11'd232;
    242: stateMap = 11'd233;
    243: stateMap = 11'd234;
    244: stateMap = 11'd235;
    245: stateMap = 11'd236;
    246: stateMap = 11'd237;
    247: stateMap = 11'd238;
    248: stateMap = 11'd239;
    249: stateMap = 11'd240;
    250: stateMap = 11'd241;
    251: stateMap = 11'd242;
    252: stateMap = 11'd243;
    253: stateMap = 11'd244;
    254: stateMap = 11'd245;
    255: stateMap = 11'd246;
    256: stateMap = 11'd247;
    257: stateMap = 11'd248;
    258: stateMap = 11'd249;
    259: stateMap = 11'd250;
    260: stateMap = 11'd251;
    261: stateMap = 11'd252;
    262: stateMap = 11'd253;
    263: stateMap = 11'd254;
    264: stateMap = 11'd255;
    265: stateMap = 11'd256;
    266: stateMap = 11'd63;
    267: stateMap = 11'd257;
    268: stateMap = 11'd258;
    269: stateMap = 11'd259;
    270: stateMap = 11'd260;
    271: stateMap = 11'd261;
    272: stateMap = 11'd246;
    273: stateMap = 11'd262;
    274: stateMap = 11'd263;
    275: stateMap = 11'd264;
    276: stateMap = 11'd265;
    277: stateMap = 11'd250;
    278: stateMap = 11'd266;
    279: stateMap = 11'd267;
    280: stateMap = 11'd268;
    281: stateMap = 11'd269;
    282: stateMap = 11'd270;
    283: stateMap = 11'd271;
    284: stateMap = 11'd272;
    285: stateMap = 11'd273;
    286: stateMap = 11'd274;
    287: stateMap = 11'd275;
    288: stateMap = 11'd276;
    289: stateMap = 11'd277;
    290: stateMap = 11'd278;
    291: stateMap = 11'd279;
    292: stateMap = 11'd280;
    293: stateMap = 11'd281;
    294: stateMap = 11'd282;
    295: stateMap = 11'd283;
    296: stateMap = 11'd284;
    297: stateMap = 11'd285;
    298: stateMap = 11'd286;
    299: stateMap = 11'd287;
    300: stateMap = 11'd288;
    301: stateMap = 11'd289;
    302: stateMap = 11'd290;
    303: stateMap = 11'd291;
    304: stateMap = 11'd292;
    305: stateMap = 11'd293;
    306: stateMap = 11'd294;
    307: stateMap = 11'd295;
    308: stateMap = 11'd296;
    309: stateMap = 11'd297;
    310: stateMap = 11'd298;
    311: stateMap = 11'd299;
    312: stateMap = 11'd300;
    313: stateMap = 11'd301;
    314: stateMap = 11'd302;
    315: stateMap = 11'd303;
    316: stateMap = 11'd304;
    317: stateMap = 11'd305;
    318: stateMap = 11'd306;
    319: stateMap = 11'd307;
    320: stateMap = 11'd308;
    321: stateMap = 11'd309;
    322: stateMap = 11'd310;
    323: stateMap = 11'd267;
    324: stateMap = 11'd311;
    325: stateMap = 11'd312;
    326: stateMap = 11'd313;
    327: stateMap = 11'd314;
    328: stateMap = 11'd315;
    329: stateMap = 11'd268;
    330: stateMap = 11'd316;
    331: stateMap = 11'd317;
    332: stateMap = 11'd249;
    333: stateMap = 11'd269;
    334: stateMap = 11'd318;
    335: stateMap = 11'd319;
    336: stateMap = 11'd320;
    337: stateMap = 11'd271;
    338: stateMap = 11'd321;
    339: stateMap = 11'd322;
    340: stateMap = 11'd323;
    341: stateMap = 11'd273;
    342: stateMap = 11'd324;
    343: stateMap = 11'd325;
    344: stateMap = 11'd326;
    345: stateMap = 11'd274;
    346: stateMap = 11'd327;
    347: stateMap = 11'd328;
    348: stateMap = 11'd329;
    349: stateMap = 11'd276;
    350: stateMap = 11'd330;
    351: stateMap = 11'd67;
    352: stateMap = 11'd331;
    353: stateMap = 11'd277;
    354: stateMap = 11'd332;
    355: stateMap = 11'd333;
    356: stateMap = 11'd334;
    357: stateMap = 11'd279;
    358: stateMap = 11'd335;
    359: stateMap = 11'd336;
    360: stateMap = 11'd337;
    361: stateMap = 11'd281;
    362: stateMap = 11'd338;
    363: stateMap = 11'd43;
    364: stateMap = 11'd339;
    365: stateMap = 11'd283;
    366: stateMap = 11'd237;
    367: stateMap = 11'd340;
    368: stateMap = 11'd341;
    369: stateMap = 11'd285;
    370: stateMap = 11'd342;
    371: stateMap = 11'd343;
    372: stateMap = 11'd287;
    373: stateMap = 11'd344;
    374: stateMap = 11'd345;
    375: stateMap = 11'd289;
    376: stateMap = 11'd291;
    377: stateMap = 11'd293;
    378: stateMap = 11'd295;
    379: stateMap = 11'd297;
    380: stateMap = 11'd298;
    381: stateMap = 11'd299;
    382: stateMap = 11'd300;
    383: stateMap = 11'd301;
    384: stateMap = 11'd302;
    385: stateMap = 11'd303;
    386: stateMap = 11'd247;
    387: stateMap = 11'd309;
    388: stateMap = 11'd346;
    389: stateMap = 11'd347;
    390: stateMap = 11'd348;
    391: stateMap = 11'd349;
    392: stateMap = 11'd348;
    393: stateMap = 11'd350;
    394: stateMap = 11'd351;
    395: stateMap = 11'd352;
    396: stateMap = 11'd353;
    397: stateMap = 11'd354;
    398: stateMap = 11'd355;
    399: stateMap = 11'd356;
    400: stateMap = 11'd357;
    401: stateMap = 11'd358;
    402: stateMap = 11'd359;
    403: stateMap = 11'd65;
    404: stateMap = 11'd359;
    405: stateMap = 11'd360;
    406: stateMap = 11'd334;
    407: stateMap = 11'd67;
    408: stateMap = 11'd352;
    409: stateMap = 11'd361;
    410: stateMap = 11'd362;
    411: stateMap = 11'd363;
    412: stateMap = 11'd364;
    413: stateMap = 11'd365;
    414: stateMap = 11'd331;
    415: stateMap = 11'd366;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b1;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b1;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b1;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b0;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b0;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b0;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b0;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b0;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b0;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b0;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b1;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b1;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b0;
    62: acceptStates = 1'b1;
    63: acceptStates = 1'b0;
    64: acceptStates = 1'b0;
    65: acceptStates = 1'b0;
    66: acceptStates = 1'b1;
    67: acceptStates = 1'b0;
    68: acceptStates = 1'b0;
    69: acceptStates = 1'b0;
    70: acceptStates = 1'b0;
    71: acceptStates = 1'b0;
    72: acceptStates = 1'b0;
    73: acceptStates = 1'b0;
    74: acceptStates = 1'b0;
    75: acceptStates = 1'b0;
    76: acceptStates = 1'b0;
    77: acceptStates = 1'b0;
    78: acceptStates = 1'b0;
    79: acceptStates = 1'b0;
    80: acceptStates = 1'b0;
    81: acceptStates = 1'b0;
    82: acceptStates = 1'b0;
    83: acceptStates = 1'b0;
    84: acceptStates = 1'b0;
    85: acceptStates = 1'b0;
    86: acceptStates = 1'b0;
    87: acceptStates = 1'b0;
    88: acceptStates = 1'b0;
    89: acceptStates = 1'b0;
    90: acceptStates = 1'b0;
    91: acceptStates = 1'b0;
    92: acceptStates = 1'b0;
    93: acceptStates = 1'b0;
    94: acceptStates = 1'b0;
    95: acceptStates = 1'b0;
    96: acceptStates = 1'b0;
    97: acceptStates = 1'b0;
    98: acceptStates = 1'b0;
    99: acceptStates = 1'b0;
    100: acceptStates = 1'b0;
    101: acceptStates = 1'b0;
    102: acceptStates = 1'b0;
    103: acceptStates = 1'b0;
    104: acceptStates = 1'b0;
    105: acceptStates = 1'b0;
    106: acceptStates = 1'b0;
    107: acceptStates = 1'b0;
    108: acceptStates = 1'b0;
    109: acceptStates = 1'b0;
    110: acceptStates = 1'b0;
    111: acceptStates = 1'b0;
    112: acceptStates = 1'b0;
    113: acceptStates = 1'b0;
    114: acceptStates = 1'b0;
    115: acceptStates = 1'b0;
    116: acceptStates = 1'b0;
    117: acceptStates = 1'b0;
    118: acceptStates = 1'b0;
    119: acceptStates = 1'b0;
    120: acceptStates = 1'b0;
    121: acceptStates = 1'b0;
    122: acceptStates = 1'b0;
    123: acceptStates = 1'b0;
    124: acceptStates = 1'b0;
    125: acceptStates = 1'b0;
    126: acceptStates = 1'b0;
    127: acceptStates = 1'b0;
    128: acceptStates = 1'b0;
    129: acceptStates = 1'b0;
    130: acceptStates = 1'b0;
    131: acceptStates = 1'b0;
    132: acceptStates = 1'b0;
    133: acceptStates = 1'b0;
    134: acceptStates = 1'b0;
    135: acceptStates = 1'b0;
    136: acceptStates = 1'b0;
    137: acceptStates = 1'b0;
    138: acceptStates = 1'b0;
    139: acceptStates = 1'b0;
    140: acceptStates = 1'b0;
    141: acceptStates = 1'b0;
    142: acceptStates = 1'b0;
    143: acceptStates = 1'b0;
    144: acceptStates = 1'b0;
    145: acceptStates = 1'b0;
    146: acceptStates = 1'b0;
    147: acceptStates = 1'b0;
    148: acceptStates = 1'b0;
    149: acceptStates = 1'b0;
    150: acceptStates = 1'b0;
    151: acceptStates = 1'b0;
    152: acceptStates = 1'b0;
    153: acceptStates = 1'b0;
    154: acceptStates = 1'b0;
    155: acceptStates = 1'b0;
    156: acceptStates = 1'b0;
    157: acceptStates = 1'b0;
    158: acceptStates = 1'b0;
    159: acceptStates = 1'b0;
    160: acceptStates = 1'b0;
    161: acceptStates = 1'b0;
    162: acceptStates = 1'b0;
    163: acceptStates = 1'b0;
    164: acceptStates = 1'b0;
    165: acceptStates = 1'b0;
    166: acceptStates = 1'b0;
    167: acceptStates = 1'b0;
    168: acceptStates = 1'b0;
    169: acceptStates = 1'b0;
    170: acceptStates = 1'b0;
    171: acceptStates = 1'b0;
    172: acceptStates = 1'b0;
    173: acceptStates = 1'b0;
    174: acceptStates = 1'b0;
    175: acceptStates = 1'b0;
    176: acceptStates = 1'b0;
    177: acceptStates = 1'b0;
    178: acceptStates = 1'b0;
    179: acceptStates = 1'b0;
    180: acceptStates = 1'b0;
    181: acceptStates = 1'b0;
    182: acceptStates = 1'b0;
    183: acceptStates = 1'b0;
    184: acceptStates = 1'b0;
    185: acceptStates = 1'b0;
    186: acceptStates = 1'b0;
    187: acceptStates = 1'b0;
    188: acceptStates = 1'b0;
    189: acceptStates = 1'b0;
    190: acceptStates = 1'b0;
    191: acceptStates = 1'b0;
    192: acceptStates = 1'b0;
    193: acceptStates = 1'b0;
    194: acceptStates = 1'b0;
    195: acceptStates = 1'b0;
    196: acceptStates = 1'b0;
    197: acceptStates = 1'b0;
    198: acceptStates = 1'b0;
    199: acceptStates = 1'b0;
    200: acceptStates = 1'b0;
    201: acceptStates = 1'b0;
    202: acceptStates = 1'b0;
    203: acceptStates = 1'b0;
    204: acceptStates = 1'b0;
    205: acceptStates = 1'b0;
    206: acceptStates = 1'b0;
    207: acceptStates = 1'b0;
    208: acceptStates = 1'b0;
    209: acceptStates = 1'b0;
    210: acceptStates = 1'b0;
    211: acceptStates = 1'b0;
    212: acceptStates = 1'b0;
    213: acceptStates = 1'b0;
    214: acceptStates = 1'b0;
    215: acceptStates = 1'b0;
    216: acceptStates = 1'b0;
    217: acceptStates = 1'b0;
    218: acceptStates = 1'b0;
    219: acceptStates = 1'b0;
    220: acceptStates = 1'b0;
    221: acceptStates = 1'b0;
    222: acceptStates = 1'b0;
    223: acceptStates = 1'b0;
    224: acceptStates = 1'b0;
    225: acceptStates = 1'b0;
    226: acceptStates = 1'b0;
    227: acceptStates = 1'b0;
    228: acceptStates = 1'b0;
    229: acceptStates = 1'b0;
    230: acceptStates = 1'b0;
    231: acceptStates = 1'b0;
    232: acceptStates = 1'b0;
    233: acceptStates = 1'b0;
    234: acceptStates = 1'b0;
    235: acceptStates = 1'b0;
    236: acceptStates = 1'b0;
    237: acceptStates = 1'b0;
    238: acceptStates = 1'b0;
    239: acceptStates = 1'b0;
    240: acceptStates = 1'b0;
    241: acceptStates = 1'b0;
    242: acceptStates = 1'b0;
    243: acceptStates = 1'b0;
    244: acceptStates = 1'b0;
    245: acceptStates = 1'b0;
    246: acceptStates = 1'b0;
    247: acceptStates = 1'b0;
    248: acceptStates = 1'b0;
    249: acceptStates = 1'b0;
    250: acceptStates = 1'b0;
    251: acceptStates = 1'b0;
    252: acceptStates = 1'b0;
    253: acceptStates = 1'b0;
    254: acceptStates = 1'b0;
    255: acceptStates = 1'b1;
    256: acceptStates = 1'b1;
    257: acceptStates = 1'b0;
    258: acceptStates = 1'b0;
    259: acceptStates = 1'b0;
    260: acceptStates = 1'b0;
    261: acceptStates = 1'b0;
    262: acceptStates = 1'b0;
    263: acceptStates = 1'b0;
    264: acceptStates = 1'b0;
    265: acceptStates = 1'b0;
    266: acceptStates = 1'b0;
    267: acceptStates = 1'b0;
    268: acceptStates = 1'b0;
    269: acceptStates = 1'b0;
    270: acceptStates = 1'b0;
    271: acceptStates = 1'b0;
    272: acceptStates = 1'b0;
    273: acceptStates = 1'b0;
    274: acceptStates = 1'b0;
    275: acceptStates = 1'b0;
    276: acceptStates = 1'b0;
    277: acceptStates = 1'b0;
    278: acceptStates = 1'b0;
    279: acceptStates = 1'b0;
    280: acceptStates = 1'b0;
    281: acceptStates = 1'b0;
    282: acceptStates = 1'b0;
    283: acceptStates = 1'b0;
    284: acceptStates = 1'b0;
    285: acceptStates = 1'b0;
    286: acceptStates = 1'b0;
    287: acceptStates = 1'b0;
    288: acceptStates = 1'b0;
    289: acceptStates = 1'b0;
    290: acceptStates = 1'b0;
    291: acceptStates = 1'b0;
    292: acceptStates = 1'b0;
    293: acceptStates = 1'b0;
    294: acceptStates = 1'b0;
    295: acceptStates = 1'b0;
    296: acceptStates = 1'b0;
    297: acceptStates = 1'b0;
    298: acceptStates = 1'b0;
    299: acceptStates = 1'b0;
    300: acceptStates = 1'b0;
    301: acceptStates = 1'b0;
    302: acceptStates = 1'b0;
    303: acceptStates = 1'b0;
    304: acceptStates = 1'b0;
    305: acceptStates = 1'b0;
    306: acceptStates = 1'b0;
    307: acceptStates = 1'b0;
    308: acceptStates = 1'b0;
    309: acceptStates = 1'b0;
    310: acceptStates = 1'b0;
    311: acceptStates = 1'b0;
    312: acceptStates = 1'b0;
    313: acceptStates = 1'b0;
    314: acceptStates = 1'b0;
    315: acceptStates = 1'b0;
    316: acceptStates = 1'b0;
    317: acceptStates = 1'b0;
    318: acceptStates = 1'b0;
    319: acceptStates = 1'b0;
    320: acceptStates = 1'b0;
    321: acceptStates = 1'b1;
    322: acceptStates = 1'b0;
    323: acceptStates = 1'b0;
    324: acceptStates = 1'b0;
    325: acceptStates = 1'b0;
    326: acceptStates = 1'b0;
    327: acceptStates = 1'b0;
    328: acceptStates = 1'b0;
    329: acceptStates = 1'b0;
    330: acceptStates = 1'b0;
    331: acceptStates = 1'b0;
    332: acceptStates = 1'b0;
    333: acceptStates = 1'b0;
    334: acceptStates = 1'b0;
    335: acceptStates = 1'b0;
    336: acceptStates = 1'b0;
    337: acceptStates = 1'b0;
    338: acceptStates = 1'b0;
    339: acceptStates = 1'b0;
    340: acceptStates = 1'b0;
    341: acceptStates = 1'b0;
    342: acceptStates = 1'b0;
    343: acceptStates = 1'b0;
    344: acceptStates = 1'b0;
    345: acceptStates = 1'b0;
    346: acceptStates = 1'b0;
    347: acceptStates = 1'b0;
    348: acceptStates = 1'b0;
    349: acceptStates = 1'b0;
    350: acceptStates = 1'b0;
    351: acceptStates = 1'b0;
    352: acceptStates = 1'b0;
    353: acceptStates = 1'b0;
    354: acceptStates = 1'b0;
    355: acceptStates = 1'b0;
    356: acceptStates = 1'b0;
    357: acceptStates = 1'b0;
    358: acceptStates = 1'b0;
    359: acceptStates = 1'b0;
    360: acceptStates = 1'b0;
    361: acceptStates = 1'b0;
    362: acceptStates = 1'b0;
    363: acceptStates = 1'b0;
    364: acceptStates = 1'b0;
    365: acceptStates = 1'b0;
    366: acceptStates = 1'b0;
    367: acceptStates = 1'b0;
    368: acceptStates = 1'b0;
    369: acceptStates = 1'b0;
    370: acceptStates = 1'b0;
    371: acceptStates = 1'b0;
    372: acceptStates = 1'b0;
    373: acceptStates = 1'b0;
    374: acceptStates = 1'b0;
    375: acceptStates = 1'b0;
    376: acceptStates = 1'b0;
    377: acceptStates = 1'b0;
    378: acceptStates = 1'b0;
    379: acceptStates = 1'b0;
    380: acceptStates = 1'b0;
    381: acceptStates = 1'b0;
    382: acceptStates = 1'b0;
    383: acceptStates = 1'b0;
    384: acceptStates = 1'b0;
    385: acceptStates = 1'b0;
    386: acceptStates = 1'b0;
    387: acceptStates = 1'b0;
    388: acceptStates = 1'b0;
    389: acceptStates = 1'b0;
    390: acceptStates = 1'b1;
    391: acceptStates = 1'b0;
    392: acceptStates = 1'b0;
    393: acceptStates = 1'b0;
    394: acceptStates = 1'b0;
    395: acceptStates = 1'b0;
    396: acceptStates = 1'b0;
    397: acceptStates = 1'b0;
    398: acceptStates = 1'b0;
    399: acceptStates = 1'b0;
    400: acceptStates = 1'b0;
    401: acceptStates = 1'b0;
    402: acceptStates = 1'b1;
    403: acceptStates = 1'b0;
    404: acceptStates = 1'b0;
    405: acceptStates = 1'b0;
    406: acceptStates = 1'b0;
    407: acceptStates = 1'b0;
    408: acceptStates = 1'b0;
    409: acceptStates = 1'b0;
    410: acceptStates = 1'b0;
    411: acceptStates = 1'b0;
    412: acceptStates = 1'b0;
    413: acceptStates = 1'b0;
    414: acceptStates = 1'b0;
    415: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd1;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd5;
      3: stateTransition = 11'd3;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd3;
      6: stateTransition = 11'd3;
      7: stateTransition = 11'd5;
      8: stateTransition = 11'd3;
      9: stateTransition = 11'd3;
      10: stateTransition = 11'd3;
      11: stateTransition = 11'd3;
      12: stateTransition = 11'd3;
      13: stateTransition = 11'd3;
      14: stateTransition = 11'd3;
      15: stateTransition = 11'd3;
      16: stateTransition = 11'd3;
      17: stateTransition = 11'd3;
      18: stateTransition = 11'd3;
      19: stateTransition = 11'd3;
      20: stateTransition = 11'd3;
      21: stateTransition = 11'd3;
      22: stateTransition = 11'd3;
      23: stateTransition = 11'd3;
      24: stateTransition = 11'd3;
      25: stateTransition = 11'd3;
      26: stateTransition = 11'd3;
      27: stateTransition = 11'd3;
      28: stateTransition = 11'd3;
      29: stateTransition = 11'd3;
      30: stateTransition = 11'd3;
      31: stateTransition = 11'd3;
      32: stateTransition = 11'd3;
      33: stateTransition = 11'd3;
      34: stateTransition = 11'd3;
      35: stateTransition = 11'd3;
      36: stateTransition = 11'd3;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd47;
      2: stateTransition = 11'd257;
      3: stateTransition = 11'd47;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd47;
      6: stateTransition = 11'd47;
      7: stateTransition = 11'd257;
      8: stateTransition = 11'd47;
      9: stateTransition = 11'd47;
      10: stateTransition = 11'd47;
      11: stateTransition = 11'd47;
      12: stateTransition = 11'd47;
      13: stateTransition = 11'd47;
      14: stateTransition = 11'd47;
      15: stateTransition = 11'd47;
      16: stateTransition = 11'd47;
      17: stateTransition = 11'd47;
      18: stateTransition = 11'd47;
      19: stateTransition = 11'd47;
      20: stateTransition = 11'd47;
      21: stateTransition = 11'd47;
      22: stateTransition = 11'd47;
      23: stateTransition = 11'd47;
      24: stateTransition = 11'd47;
      25: stateTransition = 11'd47;
      26: stateTransition = 11'd47;
      27: stateTransition = 11'd47;
      28: stateTransition = 11'd47;
      29: stateTransition = 11'd47;
      30: stateTransition = 11'd47;
      31: stateTransition = 11'd47;
      32: stateTransition = 11'd47;
      33: stateTransition = 11'd47;
      34: stateTransition = 11'd47;
      35: stateTransition = 11'd47;
      36: stateTransition = 11'd47;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd322;
      2: stateTransition = 11'd48;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd322;
      7: stateTransition = 11'd48;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd322;
      10: stateTransition = 11'd322;
      11: stateTransition = 11'd322;
      12: stateTransition = 11'd322;
      13: stateTransition = 11'd322;
      14: stateTransition = 11'd322;
      15: stateTransition = 11'd322;
      16: stateTransition = 11'd322;
      17: stateTransition = 11'd322;
      18: stateTransition = 11'd322;
      19: stateTransition = 11'd322;
      20: stateTransition = 11'd322;
      21: stateTransition = 11'd322;
      22: stateTransition = 11'd322;
      23: stateTransition = 11'd322;
      24: stateTransition = 11'd322;
      25: stateTransition = 11'd322;
      26: stateTransition = 11'd322;
      27: stateTransition = 11'd322;
      28: stateTransition = 11'd322;
      29: stateTransition = 11'd322;
      30: stateTransition = 11'd322;
      31: stateTransition = 11'd322;
      32: stateTransition = 11'd322;
      33: stateTransition = 11'd322;
      34: stateTransition = 11'd59;
      35: stateTransition = 11'd59;
      36: stateTransition = 11'd322;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd7;
      3: stateTransition = 11'd7;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd7;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd7;
      8: stateTransition = 11'd7;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd7;
      35: stateTransition = 11'd7;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd14;
      2: stateTransition = 11'd410;
      3: stateTransition = 11'd14;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd14;
      6: stateTransition = 11'd14;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd14;
      9: stateTransition = 11'd14;
      10: stateTransition = 11'd14;
      11: stateTransition = 11'd14;
      12: stateTransition = 11'd14;
      13: stateTransition = 11'd14;
      14: stateTransition = 11'd14;
      15: stateTransition = 11'd14;
      16: stateTransition = 11'd14;
      17: stateTransition = 11'd14;
      18: stateTransition = 11'd14;
      19: stateTransition = 11'd14;
      20: stateTransition = 11'd14;
      21: stateTransition = 11'd14;
      22: stateTransition = 11'd14;
      23: stateTransition = 11'd14;
      24: stateTransition = 11'd14;
      25: stateTransition = 11'd14;
      26: stateTransition = 11'd14;
      27: stateTransition = 11'd14;
      28: stateTransition = 11'd14;
      29: stateTransition = 11'd14;
      30: stateTransition = 11'd14;
      31: stateTransition = 11'd14;
      32: stateTransition = 11'd14;
      33: stateTransition = 11'd14;
      34: stateTransition = 11'd14;
      35: stateTransition = 11'd14;
      36: stateTransition = 11'd14;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd327;
      2: stateTransition = 11'd408;
      3: stateTransition = 11'd403;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd69;
      6: stateTransition = 11'd69;
      7: stateTransition = 11'd270;
      8: stateTransition = 11'd328;
      9: stateTransition = 11'd69;
      10: stateTransition = 11'd69;
      11: stateTransition = 11'd69;
      12: stateTransition = 11'd69;
      13: stateTransition = 11'd69;
      14: stateTransition = 11'd69;
      15: stateTransition = 11'd69;
      16: stateTransition = 11'd69;
      17: stateTransition = 11'd69;
      18: stateTransition = 11'd69;
      19: stateTransition = 11'd69;
      20: stateTransition = 11'd69;
      21: stateTransition = 11'd69;
      22: stateTransition = 11'd69;
      23: stateTransition = 11'd69;
      24: stateTransition = 11'd69;
      25: stateTransition = 11'd69;
      26: stateTransition = 11'd69;
      27: stateTransition = 11'd69;
      28: stateTransition = 11'd69;
      29: stateTransition = 11'd69;
      30: stateTransition = 11'd69;
      31: stateTransition = 11'd69;
      32: stateTransition = 11'd69;
      33: stateTransition = 11'd69;
      34: stateTransition = 11'd403;
      35: stateTransition = 11'd328;
      36: stateTransition = 11'd327;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd327;
      2: stateTransition = 11'd408;
      3: stateTransition = 11'd403;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd403;
      6: stateTransition = 11'd69;
      7: stateTransition = 11'd270;
      8: stateTransition = 11'd328;
      9: stateTransition = 11'd69;
      10: stateTransition = 11'd69;
      11: stateTransition = 11'd69;
      12: stateTransition = 11'd69;
      13: stateTransition = 11'd69;
      14: stateTransition = 11'd69;
      15: stateTransition = 11'd69;
      16: stateTransition = 11'd69;
      17: stateTransition = 11'd69;
      18: stateTransition = 11'd69;
      19: stateTransition = 11'd69;
      20: stateTransition = 11'd69;
      21: stateTransition = 11'd69;
      22: stateTransition = 11'd69;
      23: stateTransition = 11'd69;
      24: stateTransition = 11'd69;
      25: stateTransition = 11'd69;
      26: stateTransition = 11'd69;
      27: stateTransition = 11'd69;
      28: stateTransition = 11'd69;
      29: stateTransition = 11'd69;
      30: stateTransition = 11'd69;
      31: stateTransition = 11'd69;
      32: stateTransition = 11'd69;
      33: stateTransition = 11'd69;
      34: stateTransition = 11'd403;
      35: stateTransition = 11'd328;
      36: stateTransition = 11'd327;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd395;
      3: stateTransition = 11'd332;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd332;
      6: stateTransition = 11'd332;
      7: stateTransition = 11'd270;
      8: stateTransition = 11'd336;
      9: stateTransition = 11'd332;
      10: stateTransition = 11'd332;
      11: stateTransition = 11'd332;
      12: stateTransition = 11'd332;
      13: stateTransition = 11'd332;
      14: stateTransition = 11'd332;
      15: stateTransition = 11'd332;
      16: stateTransition = 11'd332;
      17: stateTransition = 11'd332;
      18: stateTransition = 11'd332;
      19: stateTransition = 11'd332;
      20: stateTransition = 11'd332;
      21: stateTransition = 11'd332;
      22: stateTransition = 11'd332;
      23: stateTransition = 11'd332;
      24: stateTransition = 11'd332;
      25: stateTransition = 11'd332;
      26: stateTransition = 11'd332;
      27: stateTransition = 11'd332;
      28: stateTransition = 11'd332;
      29: stateTransition = 11'd332;
      30: stateTransition = 11'd332;
      31: stateTransition = 11'd332;
      32: stateTransition = 11'd332;
      33: stateTransition = 11'd332;
      34: stateTransition = 11'd332;
      35: stateTransition = 11'd336;
      36: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd339;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd339;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd245;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd39;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd40;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd39;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd41;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd42;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd43;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd156;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd44;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd44;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd156;
      25: stateTransition = 11'd44;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd160;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd44;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd7;
      3: stateTransition = 11'd7;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd7;
      8: stateTransition = 11'd7;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd7;
      35: stateTransition = 11'd7;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd250;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd251;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd2;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd255;
      36: stateTransition = 11'd46;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd390;
      36: stateTransition = 11'd6;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd402;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd256;
      36: stateTransition = 11'd8;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd44;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd44;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd44;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd388;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd44;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd44;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd196;
      3: stateTransition = 11'd196;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd196;
      6: stateTransition = 11'd195;
      7: stateTransition = 11'd196;
      8: stateTransition = 11'd196;
      9: stateTransition = 11'd195;
      10: stateTransition = 11'd195;
      11: stateTransition = 11'd195;
      12: stateTransition = 11'd195;
      13: stateTransition = 11'd195;
      14: stateTransition = 11'd195;
      15: stateTransition = 11'd195;
      16: stateTransition = 11'd195;
      17: stateTransition = 11'd195;
      18: stateTransition = 11'd195;
      19: stateTransition = 11'd195;
      20: stateTransition = 11'd195;
      21: stateTransition = 11'd195;
      22: stateTransition = 11'd195;
      23: stateTransition = 11'd195;
      24: stateTransition = 11'd195;
      25: stateTransition = 11'd195;
      26: stateTransition = 11'd195;
      27: stateTransition = 11'd195;
      28: stateTransition = 11'd195;
      29: stateTransition = 11'd195;
      30: stateTransition = 11'd195;
      31: stateTransition = 11'd195;
      32: stateTransition = 11'd195;
      33: stateTransition = 11'd195;
      34: stateTransition = 11'd196;
      35: stateTransition = 11'd196;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd9;
      2: stateTransition = 11'd63;
      3: stateTransition = 11'd9;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd9;
      6: stateTransition = 11'd9;
      7: stateTransition = 11'd63;
      8: stateTransition = 11'd9;
      9: stateTransition = 11'd9;
      10: stateTransition = 11'd9;
      11: stateTransition = 11'd9;
      12: stateTransition = 11'd9;
      13: stateTransition = 11'd9;
      14: stateTransition = 11'd9;
      15: stateTransition = 11'd9;
      16: stateTransition = 11'd9;
      17: stateTransition = 11'd9;
      18: stateTransition = 11'd9;
      19: stateTransition = 11'd9;
      20: stateTransition = 11'd9;
      21: stateTransition = 11'd9;
      22: stateTransition = 11'd9;
      23: stateTransition = 11'd9;
      24: stateTransition = 11'd9;
      25: stateTransition = 11'd9;
      26: stateTransition = 11'd9;
      27: stateTransition = 11'd9;
      28: stateTransition = 11'd9;
      29: stateTransition = 11'd9;
      30: stateTransition = 11'd9;
      31: stateTransition = 11'd9;
      32: stateTransition = 11'd9;
      33: stateTransition = 11'd9;
      34: stateTransition = 11'd9;
      35: stateTransition = 11'd9;
      36: stateTransition = 11'd9;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd266;
      3: stateTransition = 11'd326;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd10;
      6: stateTransition = 11'd11;
      7: stateTransition = 11'd266;
      8: stateTransition = 11'd326;
      9: stateTransition = 11'd11;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd11;
      17: stateTransition = 11'd11;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd11;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      32: stateTransition = 11'd11;
      33: stateTransition = 11'd11;
      34: stateTransition = 11'd326;
      35: stateTransition = 11'd326;
      36: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd55;
      8: stateTransition = 11'd55;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd38;
      35: stateTransition = 11'd55;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd158;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd44;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd58;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd62;
      36: stateTransition = 11'd66;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd277;
      10: stateTransition = 11'd279;
      11: stateTransition = 11'd280;
      12: stateTransition = 11'd281;
      13: stateTransition = 11'd283;
      14: stateTransition = 11'd285;
      15: stateTransition = 11'd286;
      16: stateTransition = 11'd288;
      17: stateTransition = 11'd289;
      18: stateTransition = 11'd291;
      19: stateTransition = 11'd293;
      20: stateTransition = 11'd295;
      21: stateTransition = 11'd297;
      22: stateTransition = 11'd299;
      23: stateTransition = 11'd301;
      24: stateTransition = 11'd303;
      25: stateTransition = 11'd305;
      26: stateTransition = 11'd307;
      27: stateTransition = 11'd309;
      28: stateTransition = 11'd310;
      29: stateTransition = 11'd311;
      30: stateTransition = 11'd312;
      31: stateTransition = 11'd313;
      32: stateTransition = 11'd314;
      33: stateTransition = 11'd315;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd321;
      36: stateTransition = 11'd6;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd402;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd88;
      10: stateTransition = 11'd90;
      11: stateTransition = 11'd92;
      12: stateTransition = 11'd94;
      13: stateTransition = 11'd96;
      14: stateTransition = 11'd98;
      15: stateTransition = 11'd100;
      16: stateTransition = 11'd102;
      17: stateTransition = 11'd104;
      18: stateTransition = 11'd106;
      19: stateTransition = 11'd108;
      20: stateTransition = 11'd110;
      21: stateTransition = 11'd112;
      22: stateTransition = 11'd114;
      23: stateTransition = 11'd116;
      24: stateTransition = 11'd118;
      25: stateTransition = 11'd120;
      26: stateTransition = 11'd122;
      27: stateTransition = 11'd124;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd128;
      30: stateTransition = 11'd130;
      31: stateTransition = 11'd132;
      32: stateTransition = 11'd134;
      33: stateTransition = 11'd136;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd256;
      36: stateTransition = 11'd8;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd320;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd405;
      2: stateTransition = 11'd67;
      3: stateTransition = 11'd268;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd12;
      6: stateTransition = 11'd12;
      7: stateTransition = 11'd67;
      8: stateTransition = 11'd268;
      9: stateTransition = 11'd12;
      10: stateTransition = 11'd12;
      11: stateTransition = 11'd12;
      12: stateTransition = 11'd12;
      13: stateTransition = 11'd12;
      14: stateTransition = 11'd12;
      15: stateTransition = 11'd12;
      16: stateTransition = 11'd12;
      17: stateTransition = 11'd12;
      18: stateTransition = 11'd12;
      19: stateTransition = 11'd12;
      20: stateTransition = 11'd12;
      21: stateTransition = 11'd12;
      22: stateTransition = 11'd12;
      23: stateTransition = 11'd12;
      24: stateTransition = 11'd12;
      25: stateTransition = 11'd12;
      26: stateTransition = 11'd12;
      27: stateTransition = 11'd12;
      28: stateTransition = 11'd12;
      29: stateTransition = 11'd12;
      30: stateTransition = 11'd12;
      31: stateTransition = 11'd12;
      32: stateTransition = 11'd12;
      33: stateTransition = 11'd12;
      34: stateTransition = 11'd268;
      35: stateTransition = 11'd268;
      36: stateTransition = 11'd405;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd317;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd88;
      10: stateTransition = 11'd90;
      11: stateTransition = 11'd92;
      12: stateTransition = 11'd94;
      13: stateTransition = 11'd96;
      14: stateTransition = 11'd98;
      15: stateTransition = 11'd100;
      16: stateTransition = 11'd102;
      17: stateTransition = 11'd104;
      18: stateTransition = 11'd106;
      19: stateTransition = 11'd108;
      20: stateTransition = 11'd110;
      21: stateTransition = 11'd112;
      22: stateTransition = 11'd114;
      23: stateTransition = 11'd116;
      24: stateTransition = 11'd118;
      25: stateTransition = 11'd120;
      26: stateTransition = 11'd122;
      27: stateTransition = 11'd124;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd128;
      30: stateTransition = 11'd130;
      31: stateTransition = 11'd132;
      32: stateTransition = 11'd134;
      33: stateTransition = 11'd136;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    60: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd413;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd397;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd397;
      6: stateTransition = 11'd413;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd397;
      9: stateTransition = 11'd413;
      10: stateTransition = 11'd413;
      11: stateTransition = 11'd413;
      12: stateTransition = 11'd413;
      13: stateTransition = 11'd413;
      14: stateTransition = 11'd413;
      15: stateTransition = 11'd413;
      16: stateTransition = 11'd413;
      17: stateTransition = 11'd413;
      18: stateTransition = 11'd413;
      19: stateTransition = 11'd413;
      20: stateTransition = 11'd413;
      21: stateTransition = 11'd413;
      22: stateTransition = 11'd413;
      23: stateTransition = 11'd413;
      24: stateTransition = 11'd413;
      25: stateTransition = 11'd413;
      26: stateTransition = 11'd413;
      27: stateTransition = 11'd413;
      28: stateTransition = 11'd413;
      29: stateTransition = 11'd413;
      30: stateTransition = 11'd413;
      31: stateTransition = 11'd413;
      32: stateTransition = 11'd413;
      33: stateTransition = 11'd413;
      34: stateTransition = 11'd397;
      35: stateTransition = 11'd397;
      36: stateTransition = 11'd413;
      default: stateTransition = 11'bX;
    endcase
    61: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    62: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd31;
      3: stateTransition = 11'd31;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd31;
      6: stateTransition = 11'd30;
      7: stateTransition = 11'd31;
      8: stateTransition = 11'd31;
      9: stateTransition = 11'd30;
      10: stateTransition = 11'd30;
      11: stateTransition = 11'd30;
      12: stateTransition = 11'd30;
      13: stateTransition = 11'd30;
      14: stateTransition = 11'd30;
      15: stateTransition = 11'd30;
      16: stateTransition = 11'd30;
      17: stateTransition = 11'd30;
      18: stateTransition = 11'd30;
      19: stateTransition = 11'd30;
      20: stateTransition = 11'd30;
      21: stateTransition = 11'd30;
      22: stateTransition = 11'd30;
      23: stateTransition = 11'd30;
      24: stateTransition = 11'd30;
      25: stateTransition = 11'd30;
      26: stateTransition = 11'd30;
      27: stateTransition = 11'd30;
      28: stateTransition = 11'd30;
      29: stateTransition = 11'd30;
      30: stateTransition = 11'd30;
      31: stateTransition = 11'd30;
      32: stateTransition = 11'd30;
      33: stateTransition = 11'd30;
      34: stateTransition = 11'd31;
      35: stateTransition = 11'd31;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    63: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd413;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd397;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd391;
      6: stateTransition = 11'd391;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd397;
      9: stateTransition = 11'd391;
      10: stateTransition = 11'd391;
      11: stateTransition = 11'd391;
      12: stateTransition = 11'd391;
      13: stateTransition = 11'd391;
      14: stateTransition = 11'd391;
      15: stateTransition = 11'd391;
      16: stateTransition = 11'd391;
      17: stateTransition = 11'd391;
      18: stateTransition = 11'd391;
      19: stateTransition = 11'd391;
      20: stateTransition = 11'd391;
      21: stateTransition = 11'd391;
      22: stateTransition = 11'd391;
      23: stateTransition = 11'd391;
      24: stateTransition = 11'd391;
      25: stateTransition = 11'd391;
      26: stateTransition = 11'd391;
      27: stateTransition = 11'd391;
      28: stateTransition = 11'd391;
      29: stateTransition = 11'd391;
      30: stateTransition = 11'd391;
      31: stateTransition = 11'd391;
      32: stateTransition = 11'd391;
      33: stateTransition = 11'd391;
      34: stateTransition = 11'd397;
      35: stateTransition = 11'd397;
      36: stateTransition = 11'd413;
      default: stateTransition = 11'bX;
    endcase
    64: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd57;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    65: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd414;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    66: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd57;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    67: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd343;
      3: stateTransition = 11'd343;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd406;
      6: stateTransition = 11'd406;
      7: stateTransition = 11'd343;
      8: stateTransition = 11'd343;
      9: stateTransition = 11'd406;
      10: stateTransition = 11'd406;
      11: stateTransition = 11'd406;
      12: stateTransition = 11'd406;
      13: stateTransition = 11'd406;
      14: stateTransition = 11'd406;
      15: stateTransition = 11'd406;
      16: stateTransition = 11'd406;
      17: stateTransition = 11'd406;
      18: stateTransition = 11'd406;
      19: stateTransition = 11'd406;
      20: stateTransition = 11'd406;
      21: stateTransition = 11'd406;
      22: stateTransition = 11'd406;
      23: stateTransition = 11'd406;
      24: stateTransition = 11'd406;
      25: stateTransition = 11'd406;
      26: stateTransition = 11'd406;
      27: stateTransition = 11'd406;
      28: stateTransition = 11'd406;
      29: stateTransition = 11'd406;
      30: stateTransition = 11'd406;
      31: stateTransition = 11'd406;
      32: stateTransition = 11'd406;
      33: stateTransition = 11'd406;
      34: stateTransition = 11'd343;
      35: stateTransition = 11'd343;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    68: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    69: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd57;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    70: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd15;
      11: stateTransition = 11'd260;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd324;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    71: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd57;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    72: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd364;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    73: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd318;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd57;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    74: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    75: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd57;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    76: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd368;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    77: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd57;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    78: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd330;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    79: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd319;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    80: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd324;
      15: stateTransition = 11'd334;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd324;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd324;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    81: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd57;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    82: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd338;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd324;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    83: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd49;
      11: stateTransition = 11'd60;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    84: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    85: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    86: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd324;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd342;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd324;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    87: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    88: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd324;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd371;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd346;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd324;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd324;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    89: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd70;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    90: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd324;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    91: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd72;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    92: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    93: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd74;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    94: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd374;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd324;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    95: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd76;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    96: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    97: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    98: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd350;
      10: stateTransition = 11'd354;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    99: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd64;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd78;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    100: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd324;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    101: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd64;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd80;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd394;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    102: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd324;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd324;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    103: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    104: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd324;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd324;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    105: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    106: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd324;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd324;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd324;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd324;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd324;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd324;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    107: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd82;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    108: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd324;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    109: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    110: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd324;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd324;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    111: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd84;
      10: stateTransition = 11'd86;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    112: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd324;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    113: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    114: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd324;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    115: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    116: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd324;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    117: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    118: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd324;
      11: stateTransition = 11'd324;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd324;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd324;
      16: stateTransition = 11'd324;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd324;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd324;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd324;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd324;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    119: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    120: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd16;
      11: stateTransition = 11'd17;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd50;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    121: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    122: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd233;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    123: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    124: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    125: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    126: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd234;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    127: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    128: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd18;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    129: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    130: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd50;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd50;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    131: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    132: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd20;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd50;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    133: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    134: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    135: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd317;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    136: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd50;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd21;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    137: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd50;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd235;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd22;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd50;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    138: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    139: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd50;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    140: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd57;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    141: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    142: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd57;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    143: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd236;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd50;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    144: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd318;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd57;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    145: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    146: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd319;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    147: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd23;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    148: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd57;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    149: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd50;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    150: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    151: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd50;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    152: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd57;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    153: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd50;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    154: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd57;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    155: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd50;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd50;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd50;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd50;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    156: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd57;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    157: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd50;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    158: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd57;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    159: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd50;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd50;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    160: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd50;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    161: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    162: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    163: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd50;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd50;
      16: stateTransition = 11'd50;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd50;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd50;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd50;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    164: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd25;
      11: stateTransition = 11'd51;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd61;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    165: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd237;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    166: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    167: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    168: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd26;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    169: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd61;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd61;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    170: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd28;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd61;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    171: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    172: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd61;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd29;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    173: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd61;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd239;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd415;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd61;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    174: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd61;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    175: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    176: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd240;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd61;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    177: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    178: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd65;
      10: stateTransition = 11'd52;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    179: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd61;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    180: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd61;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    181: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd61;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    182: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd61;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd61;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd61;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd61;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    183: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd61;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    184: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd61;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd61;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    185: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd61;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    186: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    187: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd61;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    188: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd61;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd61;
      16: stateTransition = 11'd61;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd61;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd61;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd61;
      30: stateTransition = 11'd61;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd61;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    189: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd31;
      3: stateTransition = 11'd31;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd31;
      8: stateTransition = 11'd31;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd31;
      35: stateTransition = 11'd31;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    190: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd138;
      11: stateTransition = 11'd140;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd142;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    191: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd269;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    192: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    193: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd271;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    194: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd144;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    195: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd142;
      15: stateTransition = 11'd146;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd142;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd142;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    196: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd148;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd142;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    197: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    198: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd142;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd150;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd142;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    199: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd142;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd275;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd396;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd142;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd142;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    200: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd142;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    201: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    202: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd276;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd142;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    203: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    204: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd154;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    205: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd142;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    206: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd142;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd142;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    207: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd142;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd142;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    208: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd142;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd142;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd142;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd142;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd142;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    209: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    210: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd142;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd142;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    211: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd142;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    212: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd142;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    213: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd142;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd142;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    214: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd142;
      11: stateTransition = 11'd142;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd142;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd142;
      16: stateTransition = 11'd142;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd142;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd142;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd142;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd142;
      30: stateTransition = 11'd142;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd142;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    215: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd241;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    216: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd242;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    217: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd32;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    218: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd366;
      15: stateTransition = 11'd33;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd366;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd366;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    219: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd34;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd366;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    220: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd366;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd35;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd366;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    221: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd366;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd243;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd370;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd366;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd366;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    222: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd244;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd366;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    223: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd373;
      10: stateTransition = 11'd261;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    224: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd61;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    225: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd61;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    226: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd61;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    227: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd61;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    228: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd44;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    229: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd44;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    230: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd44;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    231: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd404;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd386;
      8: stateTransition = 11'd386;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd44;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd404;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd404;
      35: stateTransition = 11'd386;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    232: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd50;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    233: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd50;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    234: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd50;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    235: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd50;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    236: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd50;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    237: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    238: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd50;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    239: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd254;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    240: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd50;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    241: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd61;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    242: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd61;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    243: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd56;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    244: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd61;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    245: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd45;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    246: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd197;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd199;
      10: stateTransition = 11'd200;
      11: stateTransition = 11'd201;
      12: stateTransition = 11'd202;
      13: stateTransition = 11'd203;
      14: stateTransition = 11'd204;
      15: stateTransition = 11'd205;
      16: stateTransition = 11'd206;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd208;
      19: stateTransition = 11'd209;
      20: stateTransition = 11'd210;
      21: stateTransition = 11'd211;
      22: stateTransition = 11'd212;
      23: stateTransition = 11'd213;
      24: stateTransition = 11'd214;
      25: stateTransition = 11'd215;
      26: stateTransition = 11'd216;
      27: stateTransition = 11'd217;
      28: stateTransition = 11'd218;
      29: stateTransition = 11'd219;
      30: stateTransition = 11'd220;
      31: stateTransition = 11'd221;
      32: stateTransition = 11'd222;
      33: stateTransition = 11'd223;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd198;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    247: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd277;
      10: stateTransition = 11'd279;
      11: stateTransition = 11'd280;
      12: stateTransition = 11'd281;
      13: stateTransition = 11'd283;
      14: stateTransition = 11'd285;
      15: stateTransition = 11'd286;
      16: stateTransition = 11'd288;
      17: stateTransition = 11'd289;
      18: stateTransition = 11'd291;
      19: stateTransition = 11'd293;
      20: stateTransition = 11'd295;
      21: stateTransition = 11'd297;
      22: stateTransition = 11'd299;
      23: stateTransition = 11'd301;
      24: stateTransition = 11'd303;
      25: stateTransition = 11'd305;
      26: stateTransition = 11'd307;
      27: stateTransition = 11'd309;
      28: stateTransition = 11'd310;
      29: stateTransition = 11'd311;
      30: stateTransition = 11'd312;
      31: stateTransition = 11'd313;
      32: stateTransition = 11'd314;
      33: stateTransition = 11'd315;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    248: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd266;
      3: stateTransition = 11'd326;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd326;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd266;
      8: stateTransition = 11'd326;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd393;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd393;
      19: stateTransition = 11'd393;
      20: stateTransition = 11'd393;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd393;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd393;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd326;
      35: stateTransition = 11'd326;
      36: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    249: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd352;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    250: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd49;
      11: stateTransition = 11'd60;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    251: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd163;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    252: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    253: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd2;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd171;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd173;
      13: stateTransition = 11'd174;
      14: stateTransition = 11'd175;
      15: stateTransition = 11'd176;
      16: stateTransition = 11'd177;
      17: stateTransition = 11'd178;
      18: stateTransition = 11'd179;
      19: stateTransition = 11'd180;
      20: stateTransition = 11'd181;
      21: stateTransition = 11'd182;
      22: stateTransition = 11'd183;
      23: stateTransition = 11'd184;
      24: stateTransition = 11'd185;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd187;
      27: stateTransition = 11'd188;
      28: stateTransition = 11'd189;
      29: stateTransition = 11'd190;
      30: stateTransition = 11'd191;
      31: stateTransition = 11'd192;
      32: stateTransition = 11'd193;
      33: stateTransition = 11'd194;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd255;
      36: stateTransition = 11'd46;
      default: stateTransition = 11'bX;
    endcase
    254: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd321;
      36: stateTransition = 11'd6;
      default: stateTransition = 11'bX;
    endcase
    255: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd58;
      3: stateTransition = 11'd197;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd198;
      8: stateTransition = 11'd198;
      9: stateTransition = 11'd199;
      10: stateTransition = 11'd200;
      11: stateTransition = 11'd201;
      12: stateTransition = 11'd202;
      13: stateTransition = 11'd203;
      14: stateTransition = 11'd204;
      15: stateTransition = 11'd205;
      16: stateTransition = 11'd206;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd208;
      19: stateTransition = 11'd209;
      20: stateTransition = 11'd210;
      21: stateTransition = 11'd211;
      22: stateTransition = 11'd212;
      23: stateTransition = 11'd213;
      24: stateTransition = 11'd214;
      25: stateTransition = 11'd215;
      26: stateTransition = 11'd216;
      27: stateTransition = 11'd217;
      28: stateTransition = 11'd218;
      29: stateTransition = 11'd219;
      30: stateTransition = 11'd220;
      31: stateTransition = 11'd221;
      32: stateTransition = 11'd222;
      33: stateTransition = 11'd223;
      34: stateTransition = 11'd197;
      35: stateTransition = 11'd62;
      36: stateTransition = 11'd66;
      default: stateTransition = 11'bX;
    endcase
    256: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd277;
      10: stateTransition = 11'd279;
      11: stateTransition = 11'd280;
      12: stateTransition = 11'd281;
      13: stateTransition = 11'd283;
      14: stateTransition = 11'd285;
      15: stateTransition = 11'd286;
      16: stateTransition = 11'd288;
      17: stateTransition = 11'd289;
      18: stateTransition = 11'd291;
      19: stateTransition = 11'd293;
      20: stateTransition = 11'd295;
      21: stateTransition = 11'd297;
      22: stateTransition = 11'd299;
      23: stateTransition = 11'd301;
      24: stateTransition = 11'd303;
      25: stateTransition = 11'd305;
      26: stateTransition = 11'd307;
      27: stateTransition = 11'd309;
      28: stateTransition = 11'd310;
      29: stateTransition = 11'd311;
      30: stateTransition = 11'd312;
      31: stateTransition = 11'd313;
      32: stateTransition = 11'd314;
      33: stateTransition = 11'd315;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd390;
      36: stateTransition = 11'd6;
      default: stateTransition = 11'bX;
    endcase
    257: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd407;
      3: stateTransition = 11'd343;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd406;
      6: stateTransition = 11'd406;
      7: stateTransition = 11'd407;
      8: stateTransition = 11'd343;
      9: stateTransition = 11'd406;
      10: stateTransition = 11'd406;
      11: stateTransition = 11'd406;
      12: stateTransition = 11'd406;
      13: stateTransition = 11'd406;
      14: stateTransition = 11'd406;
      15: stateTransition = 11'd406;
      16: stateTransition = 11'd406;
      17: stateTransition = 11'd406;
      18: stateTransition = 11'd406;
      19: stateTransition = 11'd406;
      20: stateTransition = 11'd406;
      21: stateTransition = 11'd406;
      22: stateTransition = 11'd406;
      23: stateTransition = 11'd406;
      24: stateTransition = 11'd406;
      25: stateTransition = 11'd406;
      26: stateTransition = 11'd406;
      27: stateTransition = 11'd406;
      28: stateTransition = 11'd406;
      29: stateTransition = 11'd406;
      30: stateTransition = 11'd406;
      31: stateTransition = 11'd406;
      32: stateTransition = 11'd406;
      33: stateTransition = 11'd406;
      34: stateTransition = 11'd343;
      35: stateTransition = 11'd343;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    258: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd335;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd258;
      6: stateTransition = 11'd258;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd335;
      9: stateTransition = 11'd258;
      10: stateTransition = 11'd258;
      11: stateTransition = 11'd258;
      12: stateTransition = 11'd258;
      13: stateTransition = 11'd258;
      14: stateTransition = 11'd258;
      15: stateTransition = 11'd258;
      16: stateTransition = 11'd258;
      17: stateTransition = 11'd258;
      18: stateTransition = 11'd258;
      19: stateTransition = 11'd258;
      20: stateTransition = 11'd258;
      21: stateTransition = 11'd258;
      22: stateTransition = 11'd258;
      23: stateTransition = 11'd258;
      24: stateTransition = 11'd258;
      25: stateTransition = 11'd258;
      26: stateTransition = 11'd258;
      27: stateTransition = 11'd258;
      28: stateTransition = 11'd258;
      29: stateTransition = 11'd258;
      30: stateTransition = 11'd258;
      31: stateTransition = 11'd258;
      32: stateTransition = 11'd258;
      33: stateTransition = 11'd258;
      34: stateTransition = 11'd335;
      35: stateTransition = 11'd335;
      36: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    259: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd57;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    260: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd352;
      3: stateTransition = 11'd356;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd356;
      6: stateTransition = 11'd356;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd360;
      9: stateTransition = 11'd75;
      10: stateTransition = 11'd77;
      11: stateTransition = 11'd79;
      12: stateTransition = 11'd81;
      13: stateTransition = 11'd83;
      14: stateTransition = 11'd85;
      15: stateTransition = 11'd87;
      16: stateTransition = 11'd89;
      17: stateTransition = 11'd91;
      18: stateTransition = 11'd93;
      19: stateTransition = 11'd95;
      20: stateTransition = 11'd97;
      21: stateTransition = 11'd99;
      22: stateTransition = 11'd101;
      23: stateTransition = 11'd103;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd107;
      26: stateTransition = 11'd109;
      27: stateTransition = 11'd111;
      28: stateTransition = 11'd113;
      29: stateTransition = 11'd115;
      30: stateTransition = 11'd117;
      31: stateTransition = 11'd119;
      32: stateTransition = 11'd121;
      33: stateTransition = 11'd123;
      34: stateTransition = 11'd356;
      35: stateTransition = 11'd360;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    261: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd57;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    262: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd362;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd366;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    263: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    264: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd57;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    265: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd57;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    266: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    267: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd68;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    268: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    269: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd70;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    270: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd366;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    271: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd72;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    272: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    273: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd74;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    274: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd76;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    275: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    276: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    277: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd64;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd78;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    278: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd366;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    279: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd64;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd80;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd394;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    280: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd366;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd366;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    281: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    282: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd366;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd366;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    283: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    284: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd366;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd366;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd366;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd366;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd366;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd366;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    285: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd82;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    286: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd366;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    287: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    288: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd366;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd366;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    289: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd84;
      10: stateTransition = 11'd86;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    290: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd366;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    291: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    292: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd366;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    293: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    294: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd366;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    295: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    296: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd366;
      11: stateTransition = 11'd366;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd366;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd366;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd366;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd366;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd366;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd366;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    297: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd64;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    298: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    299: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    300: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    301: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    302: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd64;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    303: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd64;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    304: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    305: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd57;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    306: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd57;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    307: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd57;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    308: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd57;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    309: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd277;
      10: stateTransition = 11'd279;
      11: stateTransition = 11'd280;
      12: stateTransition = 11'd281;
      13: stateTransition = 11'd283;
      14: stateTransition = 11'd285;
      15: stateTransition = 11'd286;
      16: stateTransition = 11'd288;
      17: stateTransition = 11'd289;
      18: stateTransition = 11'd291;
      19: stateTransition = 11'd293;
      20: stateTransition = 11'd295;
      21: stateTransition = 11'd297;
      22: stateTransition = 11'd299;
      23: stateTransition = 11'd301;
      24: stateTransition = 11'd303;
      25: stateTransition = 11'd305;
      26: stateTransition = 11'd307;
      27: stateTransition = 11'd309;
      28: stateTransition = 11'd310;
      29: stateTransition = 11'd311;
      30: stateTransition = 11'd312;
      31: stateTransition = 11'd313;
      32: stateTransition = 11'd314;
      33: stateTransition = 11'd315;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    310: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd405;
      2: stateTransition = 11'd67;
      3: stateTransition = 11'd268;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd268;
      6: stateTransition = 11'd405;
      7: stateTransition = 11'd67;
      8: stateTransition = 11'd268;
      9: stateTransition = 11'd405;
      10: stateTransition = 11'd405;
      11: stateTransition = 11'd405;
      12: stateTransition = 11'd405;
      13: stateTransition = 11'd405;
      14: stateTransition = 11'd405;
      15: stateTransition = 11'd405;
      16: stateTransition = 11'd405;
      17: stateTransition = 11'd405;
      18: stateTransition = 11'd405;
      19: stateTransition = 11'd405;
      20: stateTransition = 11'd405;
      21: stateTransition = 11'd405;
      22: stateTransition = 11'd405;
      23: stateTransition = 11'd405;
      24: stateTransition = 11'd405;
      25: stateTransition = 11'd405;
      26: stateTransition = 11'd405;
      27: stateTransition = 11'd405;
      28: stateTransition = 11'd405;
      29: stateTransition = 11'd405;
      30: stateTransition = 11'd405;
      31: stateTransition = 11'd405;
      32: stateTransition = 11'd405;
      33: stateTransition = 11'd405;
      34: stateTransition = 11'd268;
      35: stateTransition = 11'd268;
      36: stateTransition = 11'd405;
      default: stateTransition = 11'bX;
    endcase
    311: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    312: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd4;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd259;
      10: stateTransition = 11'd323;
      11: stateTransition = 11'd329;
      12: stateTransition = 11'd333;
      13: stateTransition = 11'd337;
      14: stateTransition = 11'd341;
      15: stateTransition = 11'd345;
      16: stateTransition = 11'd349;
      17: stateTransition = 11'd353;
      18: stateTransition = 11'd357;
      19: stateTransition = 11'd361;
      20: stateTransition = 11'd365;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd372;
      23: stateTransition = 11'd375;
      24: stateTransition = 11'd376;
      25: stateTransition = 11'd377;
      26: stateTransition = 11'd378;
      27: stateTransition = 11'd379;
      28: stateTransition = 11'd380;
      29: stateTransition = 11'd381;
      30: stateTransition = 11'd382;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd384;
      33: stateTransition = 11'd385;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd390;
      36: stateTransition = 11'd6;
      default: stateTransition = 11'bX;
    endcase
    313: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd327;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd331;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd403;
      6: stateTransition = 11'd403;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd331;
      9: stateTransition = 11'd403;
      10: stateTransition = 11'd403;
      11: stateTransition = 11'd403;
      12: stateTransition = 11'd403;
      13: stateTransition = 11'd403;
      14: stateTransition = 11'd403;
      15: stateTransition = 11'd403;
      16: stateTransition = 11'd403;
      17: stateTransition = 11'd403;
      18: stateTransition = 11'd403;
      19: stateTransition = 11'd403;
      20: stateTransition = 11'd403;
      21: stateTransition = 11'd403;
      22: stateTransition = 11'd403;
      23: stateTransition = 11'd403;
      24: stateTransition = 11'd403;
      25: stateTransition = 11'd403;
      26: stateTransition = 11'd403;
      27: stateTransition = 11'd403;
      28: stateTransition = 11'd403;
      29: stateTransition = 11'd403;
      30: stateTransition = 11'd403;
      31: stateTransition = 11'd403;
      32: stateTransition = 11'd403;
      33: stateTransition = 11'd403;
      34: stateTransition = 11'd331;
      35: stateTransition = 11'd331;
      36: stateTransition = 11'd327;
      default: stateTransition = 11'bX;
    endcase
    314: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd71;
      3: stateTransition = 11'd359;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd359;
      6: stateTransition = 11'd401;
      7: stateTransition = 11'd71;
      8: stateTransition = 11'd359;
      9: stateTransition = 11'd401;
      10: stateTransition = 11'd401;
      11: stateTransition = 11'd401;
      12: stateTransition = 11'd401;
      13: stateTransition = 11'd401;
      14: stateTransition = 11'd401;
      15: stateTransition = 11'd401;
      16: stateTransition = 11'd401;
      17: stateTransition = 11'd401;
      18: stateTransition = 11'd401;
      19: stateTransition = 11'd401;
      20: stateTransition = 11'd401;
      21: stateTransition = 11'd401;
      22: stateTransition = 11'd401;
      23: stateTransition = 11'd401;
      24: stateTransition = 11'd401;
      25: stateTransition = 11'd401;
      26: stateTransition = 11'd401;
      27: stateTransition = 11'd401;
      28: stateTransition = 11'd401;
      29: stateTransition = 11'd401;
      30: stateTransition = 11'd401;
      31: stateTransition = 11'd401;
      32: stateTransition = 11'd401;
      33: stateTransition = 11'd401;
      34: stateTransition = 11'd359;
      35: stateTransition = 11'd359;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    315: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd414;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd125;
      10: stateTransition = 11'd127;
      11: stateTransition = 11'd129;
      12: stateTransition = 11'd131;
      13: stateTransition = 11'd133;
      14: stateTransition = 11'd135;
      15: stateTransition = 11'd137;
      16: stateTransition = 11'd139;
      17: stateTransition = 11'd141;
      18: stateTransition = 11'd143;
      19: stateTransition = 11'd145;
      20: stateTransition = 11'd147;
      21: stateTransition = 11'd149;
      22: stateTransition = 11'd151;
      23: stateTransition = 11'd153;
      24: stateTransition = 11'd155;
      25: stateTransition = 11'd157;
      26: stateTransition = 11'd159;
      27: stateTransition = 11'd161;
      28: stateTransition = 11'd163;
      29: stateTransition = 11'd165;
      30: stateTransition = 11'd166;
      31: stateTransition = 11'd167;
      32: stateTransition = 11'd168;
      33: stateTransition = 11'd169;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    316: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd246;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    317: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd71;
      3: stateTransition = 11'd359;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd71;
      8: stateTransition = 11'd359;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd359;
      35: stateTransition = 11'd359;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    318: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd246;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    319: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd71;
      3: stateTransition = 11'd367;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd71;
      8: stateTransition = 11'd367;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd367;
      35: stateTransition = 11'd367;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    320: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd352;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd171;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd173;
      13: stateTransition = 11'd174;
      14: stateTransition = 11'd175;
      15: stateTransition = 11'd176;
      16: stateTransition = 11'd177;
      17: stateTransition = 11'd178;
      18: stateTransition = 11'd179;
      19: stateTransition = 11'd180;
      20: stateTransition = 11'd181;
      21: stateTransition = 11'd182;
      22: stateTransition = 11'd183;
      23: stateTransition = 11'd184;
      24: stateTransition = 11'd185;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd187;
      27: stateTransition = 11'd188;
      28: stateTransition = 11'd189;
      29: stateTransition = 11'd190;
      30: stateTransition = 11'd191;
      31: stateTransition = 11'd192;
      32: stateTransition = 11'd193;
      33: stateTransition = 11'd194;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    321: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd245;
      25: stateTransition = 11'd246;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    322: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd343;
      3: stateTransition = 11'd343;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd343;
      6: stateTransition = 11'd400;
      7: stateTransition = 11'd343;
      8: stateTransition = 11'd343;
      9: stateTransition = 11'd400;
      10: stateTransition = 11'd400;
      11: stateTransition = 11'd400;
      12: stateTransition = 11'd400;
      13: stateTransition = 11'd400;
      14: stateTransition = 11'd400;
      15: stateTransition = 11'd400;
      16: stateTransition = 11'd400;
      17: stateTransition = 11'd400;
      18: stateTransition = 11'd400;
      19: stateTransition = 11'd400;
      20: stateTransition = 11'd400;
      21: stateTransition = 11'd400;
      22: stateTransition = 11'd400;
      23: stateTransition = 11'd400;
      24: stateTransition = 11'd400;
      25: stateTransition = 11'd400;
      26: stateTransition = 11'd400;
      27: stateTransition = 11'd400;
      28: stateTransition = 11'd400;
      29: stateTransition = 11'd400;
      30: stateTransition = 11'd400;
      31: stateTransition = 11'd400;
      32: stateTransition = 11'd400;
      33: stateTransition = 11'd400;
      34: stateTransition = 11'd343;
      35: stateTransition = 11'd343;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    323: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    324: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd247;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd246;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    325: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd355;
      3: stateTransition = 11'd355;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd355;
      8: stateTransition = 11'd355;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd355;
      35: stateTransition = 11'd355;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    326: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd125;
      10: stateTransition = 11'd127;
      11: stateTransition = 11'd129;
      12: stateTransition = 11'd131;
      13: stateTransition = 11'd133;
      14: stateTransition = 11'd135;
      15: stateTransition = 11'd137;
      16: stateTransition = 11'd139;
      17: stateTransition = 11'd141;
      18: stateTransition = 11'd143;
      19: stateTransition = 11'd145;
      20: stateTransition = 11'd147;
      21: stateTransition = 11'd149;
      22: stateTransition = 11'd151;
      23: stateTransition = 11'd153;
      24: stateTransition = 11'd155;
      25: stateTransition = 11'd157;
      26: stateTransition = 11'd159;
      27: stateTransition = 11'd161;
      28: stateTransition = 11'd163;
      29: stateTransition = 11'd165;
      30: stateTransition = 11'd166;
      31: stateTransition = 11'd167;
      32: stateTransition = 11'd168;
      33: stateTransition = 11'd169;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    327: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd248;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    328: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd359;
      3: stateTransition = 11'd359;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd359;
      6: stateTransition = 11'd401;
      7: stateTransition = 11'd359;
      8: stateTransition = 11'd359;
      9: stateTransition = 11'd401;
      10: stateTransition = 11'd401;
      11: stateTransition = 11'd401;
      12: stateTransition = 11'd401;
      13: stateTransition = 11'd401;
      14: stateTransition = 11'd401;
      15: stateTransition = 11'd401;
      16: stateTransition = 11'd401;
      17: stateTransition = 11'd401;
      18: stateTransition = 11'd401;
      19: stateTransition = 11'd401;
      20: stateTransition = 11'd401;
      21: stateTransition = 11'd401;
      22: stateTransition = 11'd401;
      23: stateTransition = 11'd401;
      24: stateTransition = 11'd401;
      25: stateTransition = 11'd401;
      26: stateTransition = 11'd401;
      27: stateTransition = 11'd401;
      28: stateTransition = 11'd401;
      29: stateTransition = 11'd401;
      30: stateTransition = 11'd401;
      31: stateTransition = 11'd401;
      32: stateTransition = 11'd401;
      33: stateTransition = 11'd401;
      34: stateTransition = 11'd359;
      35: stateTransition = 11'd359;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    329: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd73;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd272;
      8: stateTransition = 11'd272;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd171;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd173;
      13: stateTransition = 11'd174;
      14: stateTransition = 11'd175;
      15: stateTransition = 11'd176;
      16: stateTransition = 11'd177;
      17: stateTransition = 11'd178;
      18: stateTransition = 11'd179;
      19: stateTransition = 11'd180;
      20: stateTransition = 11'd181;
      21: stateTransition = 11'd182;
      22: stateTransition = 11'd183;
      23: stateTransition = 11'd184;
      24: stateTransition = 11'd185;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd187;
      27: stateTransition = 11'd188;
      28: stateTransition = 11'd189;
      29: stateTransition = 11'd190;
      30: stateTransition = 11'd191;
      31: stateTransition = 11'd192;
      32: stateTransition = 11'd193;
      33: stateTransition = 11'd194;
      34: stateTransition = 11'd73;
      35: stateTransition = 11'd272;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    330: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd249;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    331: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd356;
      3: stateTransition = 11'd356;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd356;
      6: stateTransition = 11'd356;
      7: stateTransition = 11'd360;
      8: stateTransition = 11'd360;
      9: stateTransition = 11'd356;
      10: stateTransition = 11'd356;
      11: stateTransition = 11'd356;
      12: stateTransition = 11'd356;
      13: stateTransition = 11'd356;
      14: stateTransition = 11'd356;
      15: stateTransition = 11'd356;
      16: stateTransition = 11'd356;
      17: stateTransition = 11'd356;
      18: stateTransition = 11'd356;
      19: stateTransition = 11'd356;
      20: stateTransition = 11'd356;
      21: stateTransition = 11'd356;
      22: stateTransition = 11'd356;
      23: stateTransition = 11'd356;
      24: stateTransition = 11'd356;
      25: stateTransition = 11'd356;
      26: stateTransition = 11'd356;
      27: stateTransition = 11'd356;
      28: stateTransition = 11'd356;
      29: stateTransition = 11'd356;
      30: stateTransition = 11'd356;
      31: stateTransition = 11'd356;
      32: stateTransition = 11'd356;
      33: stateTransition = 11'd356;
      34: stateTransition = 11'd356;
      35: stateTransition = 11'd360;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    332: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd36;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd262;
      8: stateTransition = 11'd262;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd246;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd36;
      35: stateTransition = 11'd262;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    333: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd359;
      3: stateTransition = 11'd359;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd359;
      8: stateTransition = 11'd359;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd359;
      35: stateTransition = 11'd359;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    334: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    335: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd250;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    336: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd367;
      3: stateTransition = 11'd367;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd367;
      8: stateTransition = 11'd367;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd367;
      35: stateTransition = 11'd367;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    337: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd344;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd273;
      10: stateTransition = 11'd224;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd225;
      13: stateTransition = 11'd226;
      14: stateTransition = 11'd227;
      15: stateTransition = 11'd228;
      16: stateTransition = 11'd278;
      17: stateTransition = 11'd229;
      18: stateTransition = 11'd230;
      19: stateTransition = 11'd282;
      20: stateTransition = 11'd284;
      21: stateTransition = 11'd231;
      22: stateTransition = 11'd287;
      23: stateTransition = 11'd232;
      24: stateTransition = 11'd290;
      25: stateTransition = 11'd292;
      26: stateTransition = 11'd294;
      27: stateTransition = 11'd296;
      28: stateTransition = 11'd298;
      29: stateTransition = 11'd300;
      30: stateTransition = 11'd302;
      31: stateTransition = 11'd304;
      32: stateTransition = 11'd306;
      33: stateTransition = 11'd308;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    338: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd189;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    339: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd246;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    340: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd195;
      2: stateTransition = 11'd196;
      3: stateTransition = 11'd196;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd197;
      6: stateTransition = 11'd197;
      7: stateTransition = 11'd196;
      8: stateTransition = 11'd196;
      9: stateTransition = 11'd197;
      10: stateTransition = 11'd197;
      11: stateTransition = 11'd197;
      12: stateTransition = 11'd197;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd197;
      15: stateTransition = 11'd197;
      16: stateTransition = 11'd197;
      17: stateTransition = 11'd197;
      18: stateTransition = 11'd197;
      19: stateTransition = 11'd197;
      20: stateTransition = 11'd197;
      21: stateTransition = 11'd197;
      22: stateTransition = 11'd197;
      23: stateTransition = 11'd197;
      24: stateTransition = 11'd197;
      25: stateTransition = 11'd197;
      26: stateTransition = 11'd197;
      27: stateTransition = 11'd197;
      28: stateTransition = 11'd197;
      29: stateTransition = 11'd197;
      30: stateTransition = 11'd197;
      31: stateTransition = 11'd197;
      32: stateTransition = 11'd197;
      33: stateTransition = 11'd197;
      34: stateTransition = 11'd196;
      35: stateTransition = 11'd196;
      36: stateTransition = 11'd195;
      default: stateTransition = 11'bX;
    endcase
    341: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd246;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    342: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd252;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    343: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd246;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    344: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd73;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd73;
      6: stateTransition = 11'd73;
      7: stateTransition = 11'd264;
      8: stateTransition = 11'd264;
      9: stateTransition = 11'd73;
      10: stateTransition = 11'd73;
      11: stateTransition = 11'd73;
      12: stateTransition = 11'd73;
      13: stateTransition = 11'd73;
      14: stateTransition = 11'd73;
      15: stateTransition = 11'd73;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd73;
      18: stateTransition = 11'd253;
      19: stateTransition = 11'd73;
      20: stateTransition = 11'd73;
      21: stateTransition = 11'd73;
      22: stateTransition = 11'd73;
      23: stateTransition = 11'd73;
      24: stateTransition = 11'd73;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd73;
      27: stateTransition = 11'd73;
      28: stateTransition = 11'd73;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd73;
      31: stateTransition = 11'd73;
      32: stateTransition = 11'd73;
      33: stateTransition = 11'd73;
      34: stateTransition = 11'd53;
      35: stateTransition = 11'd264;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    345: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd246;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    346: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd164;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    347: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd164;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    348: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd259;
      10: stateTransition = 11'd323;
      11: stateTransition = 11'd329;
      12: stateTransition = 11'd333;
      13: stateTransition = 11'd337;
      14: stateTransition = 11'd341;
      15: stateTransition = 11'd345;
      16: stateTransition = 11'd349;
      17: stateTransition = 11'd353;
      18: stateTransition = 11'd357;
      19: stateTransition = 11'd361;
      20: stateTransition = 11'd365;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd372;
      23: stateTransition = 11'd375;
      24: stateTransition = 11'd376;
      25: stateTransition = 11'd377;
      26: stateTransition = 11'd378;
      27: stateTransition = 11'd379;
      28: stateTransition = 11'd380;
      29: stateTransition = 11'd381;
      30: stateTransition = 11'd382;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd384;
      33: stateTransition = 11'd385;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    349: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd414;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd344;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd344;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    350: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd327;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd331;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd331;
      6: stateTransition = 11'd327;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd331;
      9: stateTransition = 11'd327;
      10: stateTransition = 11'd327;
      11: stateTransition = 11'd327;
      12: stateTransition = 11'd327;
      13: stateTransition = 11'd327;
      14: stateTransition = 11'd327;
      15: stateTransition = 11'd327;
      16: stateTransition = 11'd327;
      17: stateTransition = 11'd327;
      18: stateTransition = 11'd327;
      19: stateTransition = 11'd327;
      20: stateTransition = 11'd327;
      21: stateTransition = 11'd327;
      22: stateTransition = 11'd327;
      23: stateTransition = 11'd327;
      24: stateTransition = 11'd327;
      25: stateTransition = 11'd327;
      26: stateTransition = 11'd327;
      27: stateTransition = 11'd327;
      28: stateTransition = 11'd327;
      29: stateTransition = 11'd327;
      30: stateTransition = 11'd327;
      31: stateTransition = 11'd327;
      32: stateTransition = 11'd327;
      33: stateTransition = 11'd327;
      34: stateTransition = 11'd331;
      35: stateTransition = 11'd331;
      36: stateTransition = 11'd327;
      default: stateTransition = 11'bX;
    endcase
    351: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd325;
      8: stateTransition = 11'd325;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd412;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd325;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    352: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd352;
      3: stateTransition = 11'd356;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd356;
      6: stateTransition = 11'd356;
      7: stateTransition = 11'd398;
      8: stateTransition = 11'd360;
      9: stateTransition = 11'd356;
      10: stateTransition = 11'd356;
      11: stateTransition = 11'd356;
      12: stateTransition = 11'd356;
      13: stateTransition = 11'd356;
      14: stateTransition = 11'd356;
      15: stateTransition = 11'd356;
      16: stateTransition = 11'd356;
      17: stateTransition = 11'd356;
      18: stateTransition = 11'd356;
      19: stateTransition = 11'd356;
      20: stateTransition = 11'd356;
      21: stateTransition = 11'd356;
      22: stateTransition = 11'd356;
      23: stateTransition = 11'd356;
      24: stateTransition = 11'd356;
      25: stateTransition = 11'd356;
      26: stateTransition = 11'd356;
      27: stateTransition = 11'd356;
      28: stateTransition = 11'd356;
      29: stateTransition = 11'd356;
      30: stateTransition = 11'd356;
      31: stateTransition = 11'd356;
      32: stateTransition = 11'd356;
      33: stateTransition = 11'd356;
      34: stateTransition = 11'd356;
      35: stateTransition = 11'd360;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    353: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd37;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd265;
      8: stateTransition = 11'd265;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd412;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd37;
      35: stateTransition = 11'd265;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    354: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd351;
      3: stateTransition = 11'd355;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd411;
      6: stateTransition = 11'd411;
      7: stateTransition = 11'd351;
      8: stateTransition = 11'd355;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd411;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd411;
      20: stateTransition = 11'd411;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd355;
      35: stateTransition = 11'd355;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    355: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd356;
      3: stateTransition = 11'd356;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd356;
      6: stateTransition = 11'd356;
      7: stateTransition = 11'd360;
      8: stateTransition = 11'd360;
      9: stateTransition = 11'd75;
      10: stateTransition = 11'd77;
      11: stateTransition = 11'd79;
      12: stateTransition = 11'd81;
      13: stateTransition = 11'd83;
      14: stateTransition = 11'd85;
      15: stateTransition = 11'd87;
      16: stateTransition = 11'd89;
      17: stateTransition = 11'd91;
      18: stateTransition = 11'd93;
      19: stateTransition = 11'd95;
      20: stateTransition = 11'd97;
      21: stateTransition = 11'd99;
      22: stateTransition = 11'd101;
      23: stateTransition = 11'd103;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd107;
      26: stateTransition = 11'd109;
      27: stateTransition = 11'd111;
      28: stateTransition = 11'd113;
      29: stateTransition = 11'd115;
      30: stateTransition = 11'd117;
      31: stateTransition = 11'd119;
      32: stateTransition = 11'd121;
      33: stateTransition = 11'd123;
      34: stateTransition = 11'd356;
      35: stateTransition = 11'd360;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    356: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd71;
      3: stateTransition = 11'd367;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd367;
      6: stateTransition = 11'd363;
      7: stateTransition = 11'd71;
      8: stateTransition = 11'd367;
      9: stateTransition = 11'd363;
      10: stateTransition = 11'd363;
      11: stateTransition = 11'd363;
      12: stateTransition = 11'd363;
      13: stateTransition = 11'd363;
      14: stateTransition = 11'd363;
      15: stateTransition = 11'd363;
      16: stateTransition = 11'd363;
      17: stateTransition = 11'd363;
      18: stateTransition = 11'd363;
      19: stateTransition = 11'd363;
      20: stateTransition = 11'd363;
      21: stateTransition = 11'd363;
      22: stateTransition = 11'd363;
      23: stateTransition = 11'd363;
      24: stateTransition = 11'd363;
      25: stateTransition = 11'd363;
      26: stateTransition = 11'd363;
      27: stateTransition = 11'd363;
      28: stateTransition = 11'd363;
      29: stateTransition = 11'd363;
      30: stateTransition = 11'd363;
      31: stateTransition = 11'd363;
      32: stateTransition = 11'd363;
      33: stateTransition = 11'd363;
      34: stateTransition = 11'd367;
      35: stateTransition = 11'd367;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    357: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd355;
      3: stateTransition = 11'd355;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd355;
      6: stateTransition = 11'd347;
      7: stateTransition = 11'd355;
      8: stateTransition = 11'd355;
      9: stateTransition = 11'd347;
      10: stateTransition = 11'd347;
      11: stateTransition = 11'd347;
      12: stateTransition = 11'd347;
      13: stateTransition = 11'd347;
      14: stateTransition = 11'd347;
      15: stateTransition = 11'd347;
      16: stateTransition = 11'd347;
      17: stateTransition = 11'd347;
      18: stateTransition = 11'd347;
      19: stateTransition = 11'd347;
      20: stateTransition = 11'd347;
      21: stateTransition = 11'd347;
      22: stateTransition = 11'd347;
      23: stateTransition = 11'd347;
      24: stateTransition = 11'd347;
      25: stateTransition = 11'd347;
      26: stateTransition = 11'd347;
      27: stateTransition = 11'd347;
      28: stateTransition = 11'd347;
      29: stateTransition = 11'd347;
      30: stateTransition = 11'd347;
      31: stateTransition = 11'd347;
      32: stateTransition = 11'd347;
      33: stateTransition = 11'd347;
      34: stateTransition = 11'd355;
      35: stateTransition = 11'd355;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    358: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd363;
      2: stateTransition = 11'd367;
      3: stateTransition = 11'd367;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd367;
      6: stateTransition = 11'd363;
      7: stateTransition = 11'd367;
      8: stateTransition = 11'd367;
      9: stateTransition = 11'd363;
      10: stateTransition = 11'd363;
      11: stateTransition = 11'd363;
      12: stateTransition = 11'd363;
      13: stateTransition = 11'd363;
      14: stateTransition = 11'd363;
      15: stateTransition = 11'd363;
      16: stateTransition = 11'd363;
      17: stateTransition = 11'd363;
      18: stateTransition = 11'd363;
      19: stateTransition = 11'd363;
      20: stateTransition = 11'd363;
      21: stateTransition = 11'd363;
      22: stateTransition = 11'd363;
      23: stateTransition = 11'd363;
      24: stateTransition = 11'd363;
      25: stateTransition = 11'd363;
      26: stateTransition = 11'd363;
      27: stateTransition = 11'd363;
      28: stateTransition = 11'd363;
      29: stateTransition = 11'd363;
      30: stateTransition = 11'd363;
      31: stateTransition = 11'd363;
      32: stateTransition = 11'd363;
      33: stateTransition = 11'd363;
      34: stateTransition = 11'd367;
      35: stateTransition = 11'd367;
      36: stateTransition = 11'd363;
      default: stateTransition = 11'bX;
    endcase
    359: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    360: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd267;
      3: stateTransition = 11'd335;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd335;
      6: stateTransition = 11'd399;
      7: stateTransition = 11'd267;
      8: stateTransition = 11'd335;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd399;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd399;
      20: stateTransition = 11'd399;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd399;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd399;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd335;
      35: stateTransition = 11'd335;
      36: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    361: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd387;
      8: stateTransition = 11'd387;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd389;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd387;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    362: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd400;
      2: stateTransition = 11'd407;
      3: stateTransition = 11'd343;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd343;
      6: stateTransition = 11'd400;
      7: stateTransition = 11'd407;
      8: stateTransition = 11'd343;
      9: stateTransition = 11'd400;
      10: stateTransition = 11'd400;
      11: stateTransition = 11'd400;
      12: stateTransition = 11'd400;
      13: stateTransition = 11'd400;
      14: stateTransition = 11'd400;
      15: stateTransition = 11'd400;
      16: stateTransition = 11'd400;
      17: stateTransition = 11'd400;
      18: stateTransition = 11'd400;
      19: stateTransition = 11'd400;
      20: stateTransition = 11'd400;
      21: stateTransition = 11'd400;
      22: stateTransition = 11'd400;
      23: stateTransition = 11'd400;
      24: stateTransition = 11'd400;
      25: stateTransition = 11'd400;
      26: stateTransition = 11'd400;
      27: stateTransition = 11'd400;
      28: stateTransition = 11'd400;
      29: stateTransition = 11'd400;
      30: stateTransition = 11'd400;
      31: stateTransition = 11'd400;
      32: stateTransition = 11'd400;
      33: stateTransition = 11'd400;
      34: stateTransition = 11'd343;
      35: stateTransition = 11'd343;
      36: stateTransition = 11'd400;
      default: stateTransition = 11'bX;
    endcase
    363: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd340;
      3: stateTransition = 11'd340;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd340;
      6: stateTransition = 11'd340;
      7: stateTransition = 11'd348;
      8: stateTransition = 11'd348;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd340;
      11: stateTransition = 11'd340;
      12: stateTransition = 11'd340;
      13: stateTransition = 11'd340;
      14: stateTransition = 11'd340;
      15: stateTransition = 11'd340;
      16: stateTransition = 11'd340;
      17: stateTransition = 11'd340;
      18: stateTransition = 11'd340;
      19: stateTransition = 11'd340;
      20: stateTransition = 11'd340;
      21: stateTransition = 11'd340;
      22: stateTransition = 11'd340;
      23: stateTransition = 11'd340;
      24: stateTransition = 11'd340;
      25: stateTransition = 11'd340;
      26: stateTransition = 11'd340;
      27: stateTransition = 11'd340;
      28: stateTransition = 11'd340;
      29: stateTransition = 11'd340;
      30: stateTransition = 11'd340;
      31: stateTransition = 11'd340;
      32: stateTransition = 11'd340;
      33: stateTransition = 11'd340;
      34: stateTransition = 11'd340;
      35: stateTransition = 11'd348;
      36: stateTransition = 11'd401;
      default: stateTransition = 11'bX;
    endcase
    364: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd13;
      5: stateTransition = 11'd13;
      6: stateTransition = 11'd13;
      7: stateTransition = 11'd392;
      8: stateTransition = 11'd392;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd389;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd13;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd392;
      36: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    365: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd347;
      2: stateTransition = 11'd351;
      3: stateTransition = 11'd355;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd355;
      6: stateTransition = 11'd347;
      7: stateTransition = 11'd351;
      8: stateTransition = 11'd355;
      9: stateTransition = 11'd347;
      10: stateTransition = 11'd347;
      11: stateTransition = 11'd347;
      12: stateTransition = 11'd347;
      13: stateTransition = 11'd347;
      14: stateTransition = 11'd347;
      15: stateTransition = 11'd347;
      16: stateTransition = 11'd347;
      17: stateTransition = 11'd347;
      18: stateTransition = 11'd347;
      19: stateTransition = 11'd347;
      20: stateTransition = 11'd347;
      21: stateTransition = 11'd347;
      22: stateTransition = 11'd347;
      23: stateTransition = 11'd347;
      24: stateTransition = 11'd347;
      25: stateTransition = 11'd347;
      26: stateTransition = 11'd347;
      27: stateTransition = 11'd347;
      28: stateTransition = 11'd347;
      29: stateTransition = 11'd347;
      30: stateTransition = 11'd347;
      31: stateTransition = 11'd347;
      32: stateTransition = 11'd347;
      33: stateTransition = 11'd347;
      34: stateTransition = 11'd355;
      35: stateTransition = 11'd355;
      36: stateTransition = 11'd347;
      default: stateTransition = 11'bX;
    endcase
    366: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd30;
      2: stateTransition = 11'd263;
      3: stateTransition = 11'd404;
      4: stateTransition = 11'd37;
      5: stateTransition = 11'd404;
      6: stateTransition = 11'd404;
      7: stateTransition = 11'd54;
      8: stateTransition = 11'd54;
      9: stateTransition = 11'd404;
      10: stateTransition = 11'd404;
      11: stateTransition = 11'd404;
      12: stateTransition = 11'd404;
      13: stateTransition = 11'd404;
      14: stateTransition = 11'd404;
      15: stateTransition = 11'd404;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd404;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd404;
      20: stateTransition = 11'd404;
      21: stateTransition = 11'd404;
      22: stateTransition = 11'd404;
      23: stateTransition = 11'd404;
      24: stateTransition = 11'd404;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd404;
      27: stateTransition = 11'd409;
      28: stateTransition = 11'd404;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd404;
      31: stateTransition = 11'd404;
      32: stateTransition = 11'd404;
      33: stateTransition = 11'd404;
      34: stateTransition = 11'd263;
      35: stateTransition = 11'd54;
      36: stateTransition = 11'd30;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
