	if (fired_CATEGORY_aim) category_wd[`CATEGORY_aim] = 1 ;
	if (fired_CATEGORY_bittorrent) category_wd[`CATEGORY_bittorrent] = 1 ;
	if (fired_CATEGORY_cvs) category_wd[`CATEGORY_cvs] = 1 ;
	if (fired_CATEGORY_dhcp) category_wd[`CATEGORY_dhcp] = 1 ;
	if (fired_CATEGORY_directconnect) category_wd[`CATEGORY_directconnect] = 1 ;
	if (fired_CATEGORY_dns) category_wd[`CATEGORY_dns] = 1 ;
	if (fired_CATEGORY_fasttrack) category_wd[`CATEGORY_fasttrack] = 1 ;
	if (fired_CATEGORY_finger) category_wd[`CATEGORY_finger] = 1 ;
	if (fired_CATEGORY_freenet) category_wd[`CATEGORY_freenet] = 1 ;
	if (fired_CATEGORY_ftp) category_wd[`CATEGORY_ftp] = 1 ;
	if (fired_CATEGORY_gnutella) category_wd[`CATEGORY_gnutella] = 1 ;
	if (fired_CATEGORY_gopher) category_wd[`CATEGORY_gopher] = 1 ;
	if (fired_CATEGORY_http) category_wd[`CATEGORY_http] = 1 ;
	if (fired_CATEGORY_imap) category_wd[`CATEGORY_imap] = 1 ;
	if (fired_CATEGORY_irc) category_wd[`CATEGORY_irc] = 1 ;
	if (fired_CATEGORY_jabber) category_wd[`CATEGORY_jabber] = 1 ;
	if (fired_CATEGORY_msn) category_wd[`CATEGORY_msn] = 1 ;
	if (fired_CATEGORY_napster) category_wd[`CATEGORY_napster] = 1 ;
	if (fired_CATEGORY_netbios) category_wd[`CATEGORY_netbios] = 1 ;
	if (fired_CATEGORY_nntp) category_wd[`CATEGORY_nntp] = 1 ;
	if (fired_CATEGORY_pop3) category_wd[`CATEGORY_pop3] = 1 ;
	if (fired_CATEGORY_rlogin) category_wd[`CATEGORY_rlogin] = 1 ;
	if (fired_CATEGORY_sip) category_wd[`CATEGORY_sip] = 1 ;
	if (fired_CATEGORY_smtp) category_wd[`CATEGORY_smtp] = 1 ;
	if (fired_CATEGORY_snmp) category_wd[`CATEGORY_snmp] = 1 ;
	if (fired_CATEGORY_socks) category_wd[`CATEGORY_socks] = 1 ;
	if (fired_CATEGORY_ssh) category_wd[`CATEGORY_ssh] = 1 ;
	if (fired_CATEGORY_ssl) category_wd[`CATEGORY_ssl] = 1 ;
	if (fired_CATEGORY_subversion) category_wd[`CATEGORY_subversion] = 1 ;
	if (fired_CATEGORY_telnet) category_wd[`CATEGORY_telnet] = 1 ;
	if (fired_CATEGORY_tor) category_wd[`CATEGORY_tor] = 1 ;
	if (fired_CATEGORY_vnc) category_wd[`CATEGORY_vnc] = 1 ;
	if (fired_CATEGORY_worldofwarcraft) category_wd[`CATEGORY_worldofwarcraft] = 1 ;
	if (fired_CATEGORY_x11) category_wd[`CATEGORY_x11] = 1 ;
	if (fired_CATEGORY_yahoo) category_wd[`CATEGORY_yahoo] = 1 ;
