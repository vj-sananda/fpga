`define CATEGORY_aim 		 1
`define CATEGORY_bittorrent 		 2
`define CATEGORY_cvs 		 3
`define CATEGORY_dhcp 		 4
`define CATEGORY_directconnect 		 5
`define CATEGORY_dns 		 6
`define CATEGORY_fasttrack 		 7
`define CATEGORY_finger 		 8
`define CATEGORY_freenet 		 9
`define CATEGORY_ftp 		 10
`define CATEGORY_gnutella 		 11
`define CATEGORY_gopher 		 12
`define CATEGORY_http 		 13
`define CATEGORY_imap 		 14
`define CATEGORY_irc 		 15
`define CATEGORY_jabber 		 16
`define CATEGORY_msn 		 17
`define CATEGORY_napster 		 18
`define CATEGORY_netbios 		 19
`define CATEGORY_nntp 		 20
`define CATEGORY_pop3 		 21
`define CATEGORY_rlogin 		 22
`define CATEGORY_sip 		 23
`define CATEGORY_smtp 		 24
`define CATEGORY_snmp 		 25
`define CATEGORY_socks 		 26
`define CATEGORY_ssh 		 27
`define CATEGORY_ssl 		 28
`define CATEGORY_subversion 		 29
`define CATEGORY_telnet 		 30
`define CATEGORY_tor 		 31
`define CATEGORY_vnc 		 32
`define CATEGORY_worldofwarcraft 		 33
`define CATEGORY_x11 		 34
`define CATEGORY_yahoo 		 35
