/* ----------------------------------------------------------
 Generalized Descriptor Packer (version1: max(field_width) < input data width
 ==========================================================
 Full parameterized:
 
 Parameters: N = width of input bus
             LOG2N = ceiling( log2(M) )
             default: 8 bit ==> 32 bit ,N=8,M=4,LOG2M=2
 
 Examples: 
 
 For self test , compile this file with +define+TEST

 inputs:
   clk   => posedge triggered
   reset => active high
   din   => input data bus
   valid_din => active high, signals valid data on input bus
  
 outputs:
  
 Author: VJ Sananda
---------------------------------------------------------- */

`include "gdp.vh"

module gdp (/*AUTOARG*/
   // Outputs
   dout, valid_dout, 
   // Inputs
   clk, reset, valid_f0, valid_f1, valid_f2, valid_f3, valid_f4, 
   din_f0, din_f1, din_f2, din_f3, din_f4
   );

   parameter W = 32 ;//Width of data input bus
   parameter N = 5 ;//Number of fields in packet
   parameter LOG2N = 3 ;//Ceiling of Log2(N)
   
   parameter BIGENDIAN = 0;//1 if big endian
   
   input clk ;
   input reset ;
   
   output [W-1:0]   dout ;
   output 	   valid_dout ;

   reg [W-1:0]   dout ;
   reg 	   valid_dout ;   

   // Should be autogenerated based on packet defn
   input valid_f0 ;
   input valid_f1 ;
   input valid_f2 ;
   input valid_f3 ;
   input valid_f4 ;

   input [`F0_W-1:0] din_f0 ;
   input [`F1_W-1:0] din_f1 ;
   input [`F2_W-1:0] din_f2 ;
   input [`F3_W-1:0] din_f3 ;
   input [`F4_W-1:0] din_f4 ;

   wire valid_f0 ;
   wire valid_f1 ;
   wire valid_f2 ;
   wire valid_f3 ;
   wire valid_f4 ;

   wire [`F0_W-1:0] din_f0 ;
   wire [`F1_W-1:0] din_f1 ;
   wire [`F2_W-1:0] din_f2 ;
   wire [`F3_W-1:0] din_f3 ;
   wire [`F4_W-1:0] din_f4 ;   

   // ---------- END INPUT/OUTPUT DECL ----------

   //---------------------------------------------
   //A note about the suffixes
   //
   //   _[r,w].[c,d].[#] : choose 1 of the letters in each [] and
   //                      concatenate to build suffix
   //
   //[r,w]: r=>register, w=>wire
   //
   //[c,d]: c=>control,  d=>datapath
   //
   //[#] : Number, reflects register stage number
   //Within a clocked always block, signal on the LHS
   //of a non-blocking assignment, will have this number incremented
   //beyond the largest # of the expression on the RHS or that in a
   //conditional expression controlling the assignment
   //
   //On a wire assign, this number will not increment.
   //Goal is to make the clock cycle dependencies obvious
   //---------------------------------------------

   reg [W-1:0]	   hold_rd1 ;

   //State vector
   reg [LOG2N-1:0]   svec ;
   
   always @(posedge clk or posedge reset)
     if ( reset )
       begin
	  svec <= 0;
	  dout <= 0;
	  valid_dout <= 0;	  
       end
     else
       begin
	  valid_dout <= 0;
	  
	  case(svec)
	    0:if (valid_f0 & valid_f1 )
	      begin
		 dout[`f0_W0_MSB:`f0_W0_LSB] <= din_f0 ;
		 dout[`f1_W0_MSB:`f1_W0_LSB] <= din_f1 ;		 
		 svec <= 2 ;
	      end

	    1://if (valid_f1)
	      begin
		 svec <= 1 ;
	      end

	    2:if (valid_f2)
	      begin
		 {hold_rd1[`f2_W1_MSB:`f2_W1_LSB],dout[`f2_W0_MSB:`f2_W0_LSB]} <= din_f2 ;
		 svec <= 3 ;
		 valid_dout <= 1;
	      end

	    3:if (valid_f3)
	      begin
		 dout[`f2_W1_MSB:`f2_W1_LSB] <= hold_rd1[`f2_W1_MSB:`f2_W1_LSB] ;
		 {hold_rd1[`f3_W2_MSB:`f3_W2_LSB],dout[`f3_W1_MSB:`f3_W1_LSB]} <= din_f3 ;
		 svec <= 4 ;
		 valid_dout <= 1;
	      end

	    4:if (valid_f4)
	      begin
		 dout[`f3_W2_MSB:`f3_W2_LSB] <= hold_rd1[`f3_W2_MSB:`f3_W2_LSB] ;
		 dout[`f4_W2_MSB:`f4_W2_LSB] <= din_f4 ;		 
		 svec <= 0 ;
		 valid_dout <= 1 ;
	      end	    
	  endcase // case(svec)
       end
   
endmodule // gdp

`ifdef TEST
module test ;

   parameter W = 32 ;//Width of data input bus
   parameter N = 3 ;//Number of data words in packet
   parameter LOG2N = 2 ;//Ceiling of Log2(N)
   
   parameter BIGENDIAN = 0;//1 if big endian

   /*AUTOREGINPUT*/
   // Beginning of automatic reg inputs (for undeclared instantiated-module inputs)
   reg			clk;			// To dut of gdp.v
   reg [`F0_W-1:0]	din_f0;			// To dut of gdp.v
   reg [`F1_W-1:0]	din_f1;			// To dut of gdp.v
   reg [`F2_W-1:0]	din_f2;			// To dut of gdp.v
   reg [`F3_W-1:0]	din_f3;			// To dut of gdp.v
   reg [`F4_W-1:0]	din_f4;			// To dut of gdp.v
   reg			reset;			// To dut of gdp.v
   reg			valid_f0;		// To dut of gdp.v
   reg			valid_f1;		// To dut of gdp.v
   reg			valid_f2;		// To dut of gdp.v
   reg			valid_f3;		// To dut of gdp.v
   reg			valid_f4;		// To dut of gdp.v
   // End of automatics

   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire [W-1:0]		dout;			// From dut of gdp.v
   wire			valid_dout;		// From dut of gdp.v
   // End of automatics
   
   initial
     begin
	$dumpvars;
	clk = 0;
	din = 0;
	eop = 0;
	sop = 0;
	reset = 0;
	valid_din = 0;
	reset_dut;
	repeat(20) $display("random no = %d",$random);
       	repeat (20000) @(posedge clk);
	$finish;
     end

   always #5 clk = ~clk ;

   task reset_dut;
     begin
	@(posedge clk);
	reset <= 1;
	repeat (20) @(posedge clk);
	reset <= 0;
	repeat (20) @(posedge clk);	
     end
   endtask // reset_dut

   always @(posedge clk)
     begin
	if ($random % 4)
	  begin
	     din <= din + 1;
	     valid_din <= 1;
	  end
	else
	  valid_din <= 0;
     end

   gdp dut (/*AUTOINST*/
	    // Outputs
	    .dout			(dout[W-1:0]),
	    .valid_dout			(valid_dout),
	    // Inputs
	    .clk			(clk),
	    .reset			(reset),
	    .valid_f0			(valid_f0),
	    .valid_f1			(valid_f1),
	    .valid_f2			(valid_f2),
	    .valid_f3			(valid_f3),
	    .valid_f4			(valid_f4),
	    .din_f0			(din_f0[`F0_W-1:0]),
	    .din_f1			(din_f1[`F1_W-1:0]),
	    .din_f2			(din_f2[`F2_W-1:0]),
	    .din_f3			(din_f3[`F3_W-1:0]),
	    .din_f4			(din_f4[`F4_W-1:0]));
   

endmodule  // test

`endif

