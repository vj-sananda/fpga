`timescale 1ns/1ps

`define ENABLED_REGEX_CATEGORY_gnutella TRUE

module CATEGORY_gnutella_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_CATEGORY_gnutella

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd5;
    1: charMap = 8'd6;
    2: charMap = 8'd4;
    3: charMap = 8'd5;
    4: charMap = 8'd5;
    5: charMap = 8'd5;
    6: charMap = 8'd5;
    7: charMap = 8'd5;
    8: charMap = 8'd5;
    9: charMap = 8'd30;
    10: charMap = 8'd20;
    11: charMap = 8'd30;
    12: charMap = 8'd30;
    13: charMap = 8'd19;
    14: charMap = 8'd5;
    15: charMap = 8'd5;
    16: charMap = 8'd5;
    17: charMap = 8'd5;
    18: charMap = 8'd5;
    19: charMap = 8'd5;
    20: charMap = 8'd5;
    21: charMap = 8'd5;
    22: charMap = 8'd5;
    23: charMap = 8'd5;
    24: charMap = 8'd5;
    25: charMap = 8'd5;
    26: charMap = 8'd5;
    27: charMap = 8'd5;
    28: charMap = 8'd5;
    29: charMap = 8'd5;
    30: charMap = 8'd5;
    31: charMap = 8'd5;
    32: charMap = 8'd12;
    33: charMap = 8'd30;
    34: charMap = 8'd30;
    35: charMap = 8'd30;
    36: charMap = 8'd30;
    37: charMap = 8'd30;
    38: charMap = 8'd30;
    39: charMap = 8'd30;
    40: charMap = 8'd30;
    41: charMap = 8'd30;
    42: charMap = 8'd30;
    43: charMap = 8'd30;
    44: charMap = 8'd30;
    45: charMap = 8'd23;
    46: charMap = 8'd17;
    47: charMap = 8'd15;
    48: charMap = 8'd16;
    49: charMap = 8'd29;
    50: charMap = 8'd25;
    51: charMap = 8'd18;
    52: charMap = 8'd18;
    53: charMap = 8'd18;
    54: charMap = 8'd18;
    55: charMap = 8'd18;
    56: charMap = 8'd18;
    57: charMap = 8'd18;
    58: charMap = 8'd27;
    59: charMap = 8'd30;
    60: charMap = 8'd30;
    61: charMap = 8'd30;
    62: charMap = 8'd30;
    63: charMap = 8'd26;
    64: charMap = 8'd30;
    65: charMap = 8'd30;
    66: charMap = 8'd30;
    67: charMap = 8'd30;
    68: charMap = 8'd30;
    69: charMap = 8'd30;
    70: charMap = 8'd30;
    71: charMap = 8'd30;
    72: charMap = 8'd30;
    73: charMap = 8'd30;
    74: charMap = 8'd30;
    75: charMap = 8'd30;
    76: charMap = 8'd30;
    77: charMap = 8'd30;
    78: charMap = 8'd30;
    79: charMap = 8'd30;
    80: charMap = 8'd30;
    81: charMap = 8'd30;
    82: charMap = 8'd30;
    83: charMap = 8'd30;
    84: charMap = 8'd30;
    85: charMap = 8'd30;
    86: charMap = 8'd30;
    87: charMap = 8'd30;
    88: charMap = 8'd30;
    89: charMap = 8'd30;
    90: charMap = 8'd30;
    91: charMap = 8'd30;
    92: charMap = 8'd30;
    93: charMap = 8'd30;
    94: charMap = 8'd30;
    95: charMap = 8'd30;
    96: charMap = 8'd30;
    97: charMap = 8'd11;
    98: charMap = 8'd32;
    99: charMap = 8'd13;
    100: charMap = 8'd3;
    101: charMap = 8'd9;
    102: charMap = 8'd39;
    103: charMap = 8'd1;
    104: charMap = 8'd28;
    105: charMap = 8'd22;
    106: charMap = 8'd30;
    107: charMap = 8'd31;
    108: charMap = 8'd10;
    109: charMap = 8'd33;
    110: charMap = 8'd2;
    111: charMap = 8'd14;
    112: charMap = 8'd36;
    113: charMap = 8'd40;
    114: charMap = 8'd21;
    115: charMap = 8'd24;
    116: charMap = 8'd8;
    117: charMap = 8'd7;
    118: charMap = 8'd38;
    119: charMap = 8'd34;
    120: charMap = 8'd37;
    121: charMap = 8'd35;
    122: charMap = 8'd30;
    123: charMap = 8'd30;
    124: charMap = 8'd30;
    125: charMap = 8'd30;
    126: charMap = 8'd30;
    127: charMap = 8'd5;
    128: charMap = 8'd5;
    129: charMap = 8'd5;
    130: charMap = 8'd5;
    131: charMap = 8'd5;
    132: charMap = 8'd5;
    133: charMap = 8'd5;
    134: charMap = 8'd5;
    135: charMap = 8'd5;
    136: charMap = 8'd5;
    137: charMap = 8'd5;
    138: charMap = 8'd5;
    139: charMap = 8'd5;
    140: charMap = 8'd5;
    141: charMap = 8'd5;
    142: charMap = 8'd5;
    143: charMap = 8'd5;
    144: charMap = 8'd5;
    145: charMap = 8'd5;
    146: charMap = 8'd5;
    147: charMap = 8'd5;
    148: charMap = 8'd5;
    149: charMap = 8'd5;
    150: charMap = 8'd5;
    151: charMap = 8'd5;
    152: charMap = 8'd5;
    153: charMap = 8'd5;
    154: charMap = 8'd5;
    155: charMap = 8'd5;
    156: charMap = 8'd5;
    157: charMap = 8'd5;
    158: charMap = 8'd5;
    159: charMap = 8'd5;
    160: charMap = 8'd5;
    161: charMap = 8'd5;
    162: charMap = 8'd5;
    163: charMap = 8'd5;
    164: charMap = 8'd5;
    165: charMap = 8'd5;
    166: charMap = 8'd5;
    167: charMap = 8'd5;
    168: charMap = 8'd5;
    169: charMap = 8'd5;
    170: charMap = 8'd5;
    171: charMap = 8'd5;
    172: charMap = 8'd5;
    173: charMap = 8'd5;
    174: charMap = 8'd5;
    175: charMap = 8'd5;
    176: charMap = 8'd5;
    177: charMap = 8'd5;
    178: charMap = 8'd5;
    179: charMap = 8'd5;
    180: charMap = 8'd5;
    181: charMap = 8'd5;
    182: charMap = 8'd5;
    183: charMap = 8'd5;
    184: charMap = 8'd5;
    185: charMap = 8'd5;
    186: charMap = 8'd5;
    187: charMap = 8'd5;
    188: charMap = 8'd5;
    189: charMap = 8'd5;
    190: charMap = 8'd5;
    191: charMap = 8'd5;
    192: charMap = 8'd5;
    193: charMap = 8'd5;
    194: charMap = 8'd5;
    195: charMap = 8'd5;
    196: charMap = 8'd5;
    197: charMap = 8'd5;
    198: charMap = 8'd5;
    199: charMap = 8'd5;
    200: charMap = 8'd5;
    201: charMap = 8'd5;
    202: charMap = 8'd5;
    203: charMap = 8'd5;
    204: charMap = 8'd5;
    205: charMap = 8'd5;
    206: charMap = 8'd5;
    207: charMap = 8'd5;
    208: charMap = 8'd5;
    209: charMap = 8'd5;
    210: charMap = 8'd5;
    211: charMap = 8'd5;
    212: charMap = 8'd5;
    213: charMap = 8'd5;
    214: charMap = 8'd5;
    215: charMap = 8'd5;
    216: charMap = 8'd5;
    217: charMap = 8'd5;
    218: charMap = 8'd5;
    219: charMap = 8'd5;
    220: charMap = 8'd5;
    221: charMap = 8'd5;
    222: charMap = 8'd5;
    223: charMap = 8'd5;
    224: charMap = 8'd5;
    225: charMap = 8'd5;
    226: charMap = 8'd5;
    227: charMap = 8'd5;
    228: charMap = 8'd5;
    229: charMap = 8'd5;
    230: charMap = 8'd5;
    231: charMap = 8'd5;
    232: charMap = 8'd5;
    233: charMap = 8'd5;
    234: charMap = 8'd5;
    235: charMap = 8'd5;
    236: charMap = 8'd5;
    237: charMap = 8'd5;
    238: charMap = 8'd5;
    239: charMap = 8'd5;
    240: charMap = 8'd5;
    241: charMap = 8'd5;
    242: charMap = 8'd5;
    243: charMap = 8'd5;
    244: charMap = 8'd5;
    245: charMap = 8'd5;
    246: charMap = 8'd5;
    247: charMap = 8'd5;
    248: charMap = 8'd5;
    249: charMap = 8'd5;
    250: charMap = 8'd5;
    251: charMap = 8'd5;
    252: charMap = 8'd5;
    253: charMap = 8'd5;
    254: charMap = 8'd5;
    255: charMap = 8'd5;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd2;
    3: stateMap = 11'd3;
    4: stateMap = 11'd4;
    5: stateMap = 11'd5;
    6: stateMap = 11'd6;
    7: stateMap = 11'd7;
    8: stateMap = 11'd8;
    9: stateMap = 11'd9;
    10: stateMap = 11'd10;
    11: stateMap = 11'd11;
    12: stateMap = 11'd12;
    13: stateMap = 11'd13;
    14: stateMap = 11'd14;
    15: stateMap = 11'd15;
    16: stateMap = 11'd1;
    17: stateMap = 11'd16;
    18: stateMap = 11'd17;
    19: stateMap = 11'd18;
    20: stateMap = 11'd19;
    21: stateMap = 11'd20;
    22: stateMap = 11'd21;
    23: stateMap = 11'd22;
    24: stateMap = 11'd23;
    25: stateMap = 11'd24;
    26: stateMap = 11'd25;
    27: stateMap = 11'd12;
    28: stateMap = 11'd26;
    29: stateMap = 11'd27;
    30: stateMap = 11'd28;
    31: stateMap = 11'd29;
    32: stateMap = 11'd30;
    33: stateMap = 11'd31;
    34: stateMap = 11'd32;
    35: stateMap = 11'd33;
    36: stateMap = 11'd34;
    37: stateMap = 11'd35;
    38: stateMap = 11'd36;
    39: stateMap = 11'd37;
    40: stateMap = 11'd38;
    41: stateMap = 11'd39;
    42: stateMap = 11'd40;
    43: stateMap = 11'd41;
    44: stateMap = 11'd42;
    45: stateMap = 11'd43;
    46: stateMap = 11'd44;
    47: stateMap = 11'd45;
    48: stateMap = 11'd46;
    49: stateMap = 11'd47;
    50: stateMap = 11'd48;
    51: stateMap = 11'd49;
    52: stateMap = 11'd50;
    53: stateMap = 11'd51;
    54: stateMap = 11'd52;
    55: stateMap = 11'd53;
    56: stateMap = 11'd54;
    57: stateMap = 11'd55;
    58: stateMap = 11'd56;
    59: stateMap = 11'd57;
    60: stateMap = 11'd58;
    61: stateMap = 11'd7;
    62: stateMap = 11'd59;
    63: stateMap = 11'd60;
    64: stateMap = 11'd61;
    65: stateMap = 11'd62;
    66: stateMap = 11'd63;
    67: stateMap = 11'd64;
    68: stateMap = 11'd65;
    69: stateMap = 11'd66;
    70: stateMap = 11'd67;
    71: stateMap = 11'd68;
    72: stateMap = 11'd69;
    73: stateMap = 11'd70;
    74: stateMap = 11'd71;
    75: stateMap = 11'd72;
    76: stateMap = 11'd73;
    77: stateMap = 11'd74;
    78: stateMap = 11'd75;
    79: stateMap = 11'd2;
    80: stateMap = 11'd76;
    81: stateMap = 11'd77;
    82: stateMap = 11'd78;
    83: stateMap = 11'd79;
    84: stateMap = 11'd80;
    85: stateMap = 11'd81;
    86: stateMap = 11'd82;
    87: stateMap = 11'd83;
    88: stateMap = 11'd84;
    89: stateMap = 11'd85;
    90: stateMap = 11'd86;
    91: stateMap = 11'd87;
    92: stateMap = 11'd88;
    93: stateMap = 11'd89;
    94: stateMap = 11'd90;
    95: stateMap = 11'd91;
    96: stateMap = 11'd92;
    97: stateMap = 11'd93;
    98: stateMap = 11'd94;
    99: stateMap = 11'd95;
    100: stateMap = 11'd96;
    101: stateMap = 11'd97;
    102: stateMap = 11'd98;
    103: stateMap = 11'd99;
    104: stateMap = 11'd100;
    105: stateMap = 11'd8;
    106: stateMap = 11'd101;
    107: stateMap = 11'd102;
    108: stateMap = 11'd103;
    109: stateMap = 11'd104;
    110: stateMap = 11'd105;
    111: stateMap = 11'd106;
    112: stateMap = 11'd107;
    113: stateMap = 11'd108;
    114: stateMap = 11'd109;
    115: stateMap = 11'd110;
    116: stateMap = 11'd111;
    117: stateMap = 11'd112;
    118: stateMap = 11'd113;
    119: stateMap = 11'd114;
    120: stateMap = 11'd115;
    121: stateMap = 11'd116;
    122: stateMap = 11'd117;
    123: stateMap = 11'd118;
    124: stateMap = 11'd119;
    125: stateMap = 11'd120;
    126: stateMap = 11'd121;
    127: stateMap = 11'd122;
    128: stateMap = 11'd123;
    129: stateMap = 11'd124;
    130: stateMap = 11'd125;
    131: stateMap = 11'd126;
    132: stateMap = 11'd127;
    133: stateMap = 11'd128;
    134: stateMap = 11'd129;
    135: stateMap = 11'd130;
    136: stateMap = 11'd131;
    137: stateMap = 11'd132;
    138: stateMap = 11'd133;
    139: stateMap = 11'd134;
    140: stateMap = 11'd135;
    141: stateMap = 11'd136;
    142: stateMap = 11'd137;
    143: stateMap = 11'd138;
    144: stateMap = 11'd139;
    145: stateMap = 11'd140;
    146: stateMap = 11'd141;
    147: stateMap = 11'd142;
    148: stateMap = 11'd143;
    149: stateMap = 11'd144;
    150: stateMap = 11'd145;
    151: stateMap = 11'd146;
    152: stateMap = 11'd120;
    153: stateMap = 11'd147;
    154: stateMap = 11'd148;
    155: stateMap = 11'd149;
    156: stateMap = 11'd150;
    157: stateMap = 11'd151;
    158: stateMap = 11'd152;
    159: stateMap = 11'd153;
    160: stateMap = 11'd154;
    161: stateMap = 11'd155;
    162: stateMap = 11'd156;
    163: stateMap = 11'd157;
    164: stateMap = 11'd158;
    165: stateMap = 11'd159;
    166: stateMap = 11'd160;
    167: stateMap = 11'd161;
    168: stateMap = 11'd162;
    169: stateMap = 11'd163;
    170: stateMap = 11'd164;
    171: stateMap = 11'd165;
    172: stateMap = 11'd166;
    173: stateMap = 11'd167;
    174: stateMap = 11'd168;
    175: stateMap = 11'd169;
    176: stateMap = 11'd170;
    177: stateMap = 11'd171;
    178: stateMap = 11'd172;
    179: stateMap = 11'd173;
    180: stateMap = 11'd174;
    181: stateMap = 11'd175;
    182: stateMap = 11'd176;
    183: stateMap = 11'd177;
    184: stateMap = 11'd178;
    185: stateMap = 11'd179;
    186: stateMap = 11'd163;
    187: stateMap = 11'd180;
    188: stateMap = 11'd181;
    189: stateMap = 11'd182;
    190: stateMap = 11'd183;
    191: stateMap = 11'd125;
    192: stateMap = 11'd184;
    193: stateMap = 11'd185;
    194: stateMap = 11'd186;
    195: stateMap = 11'd187;
    196: stateMap = 11'd188;
    197: stateMap = 11'd189;
    198: stateMap = 11'd190;
    199: stateMap = 11'd191;
    200: stateMap = 11'd192;
    201: stateMap = 11'd193;
    202: stateMap = 11'd194;
    203: stateMap = 11'd195;
    204: stateMap = 11'd196;
    205: stateMap = 11'd197;
    206: stateMap = 11'd198;
    207: stateMap = 11'd199;
    208: stateMap = 11'd200;
    209: stateMap = 11'd201;
    210: stateMap = 11'd202;
    211: stateMap = 11'd203;
    212: stateMap = 11'd204;
    213: stateMap = 11'd205;
    214: stateMap = 11'd206;
    215: stateMap = 11'd207;
    216: stateMap = 11'd208;
    217: stateMap = 11'd209;
    218: stateMap = 11'd210;
    219: stateMap = 11'd211;
    220: stateMap = 11'd212;
    221: stateMap = 11'd213;
    222: stateMap = 11'd214;
    223: stateMap = 11'd215;
    224: stateMap = 11'd216;
    225: stateMap = 11'd217;
    226: stateMap = 11'd218;
    227: stateMap = 11'd219;
    228: stateMap = 11'd220;
    229: stateMap = 11'd221;
    230: stateMap = 11'd222;
    231: stateMap = 11'd223;
    232: stateMap = 11'd224;
    233: stateMap = 11'd225;
    234: stateMap = 11'd226;
    235: stateMap = 11'd227;
    236: stateMap = 11'd228;
    237: stateMap = 11'd229;
    238: stateMap = 11'd198;
    239: stateMap = 11'd230;
    240: stateMap = 11'd231;
    241: stateMap = 11'd232;
    242: stateMap = 11'd233;
    243: stateMap = 11'd234;
    244: stateMap = 11'd235;
    245: stateMap = 11'd236;
    246: stateMap = 11'd237;
    247: stateMap = 11'd238;
    248: stateMap = 11'd239;
    249: stateMap = 11'd240;
    250: stateMap = 11'd241;
    251: stateMap = 11'd242;
    252: stateMap = 11'd243;
    253: stateMap = 11'd244;
    254: stateMap = 11'd245;
    255: stateMap = 11'd246;
    256: stateMap = 11'd247;
    257: stateMap = 11'd248;
    258: stateMap = 11'd249;
    259: stateMap = 11'd250;
    260: stateMap = 11'd251;
    261: stateMap = 11'd252;
    262: stateMap = 11'd253;
    263: stateMap = 11'd254;
    264: stateMap = 11'd255;
    265: stateMap = 11'd256;
    266: stateMap = 11'd257;
    267: stateMap = 11'd258;
    268: stateMap = 11'd259;
    269: stateMap = 11'd260;
    270: stateMap = 11'd261;
    271: stateMap = 11'd262;
    272: stateMap = 11'd263;
    273: stateMap = 11'd264;
    274: stateMap = 11'd242;
    275: stateMap = 11'd265;
    276: stateMap = 11'd266;
    277: stateMap = 11'd267;
    278: stateMap = 11'd268;
    279: stateMap = 11'd269;
    280: stateMap = 11'd270;
    281: stateMap = 11'd271;
    282: stateMap = 11'd272;
    283: stateMap = 11'd273;
    284: stateMap = 11'd274;
    285: stateMap = 11'd275;
    286: stateMap = 11'd276;
    287: stateMap = 11'd277;
    288: stateMap = 11'd278;
    289: stateMap = 11'd279;
    290: stateMap = 11'd280;
    291: stateMap = 11'd281;
    292: stateMap = 11'd282;
    293: stateMap = 11'd283;
    294: stateMap = 11'd284;
    295: stateMap = 11'd285;
    296: stateMap = 11'd286;
    297: stateMap = 11'd287;
    298: stateMap = 11'd288;
    299: stateMap = 11'd289;
    300: stateMap = 11'd290;
    301: stateMap = 11'd291;
    302: stateMap = 11'd292;
    303: stateMap = 11'd293;
    304: stateMap = 11'd294;
    305: stateMap = 11'd295;
    306: stateMap = 11'd296;
    307: stateMap = 11'd297;
    308: stateMap = 11'd298;
    309: stateMap = 11'd299;
    310: stateMap = 11'd300;
    311: stateMap = 11'd301;
    312: stateMap = 11'd302;
    313: stateMap = 11'd303;
    314: stateMap = 11'd304;
    315: stateMap = 11'd305;
    316: stateMap = 11'd281;
    317: stateMap = 11'd306;
    318: stateMap = 11'd307;
    319: stateMap = 11'd308;
    320: stateMap = 11'd309;
    321: stateMap = 11'd310;
    322: stateMap = 11'd311;
    323: stateMap = 11'd312;
    324: stateMap = 11'd313;
    325: stateMap = 11'd314;
    326: stateMap = 11'd315;
    327: stateMap = 11'd316;
    328: stateMap = 11'd317;
    329: stateMap = 11'd318;
    330: stateMap = 11'd319;
    331: stateMap = 11'd320;
    332: stateMap = 11'd321;
    333: stateMap = 11'd322;
    334: stateMap = 11'd323;
    335: stateMap = 11'd324;
    336: stateMap = 11'd325;
    337: stateMap = 11'd326;
    338: stateMap = 11'd327;
    339: stateMap = 11'd328;
    340: stateMap = 11'd329;
    341: stateMap = 11'd330;
    342: stateMap = 11'd331;
    343: stateMap = 11'd332;
    344: stateMap = 11'd333;
    345: stateMap = 11'd334;
    346: stateMap = 11'd335;
    347: stateMap = 11'd336;
    348: stateMap = 11'd337;
    349: stateMap = 11'd338;
    350: stateMap = 11'd339;
    351: stateMap = 11'd340;
    352: stateMap = 11'd341;
    353: stateMap = 11'd342;
    354: stateMap = 11'd343;
    355: stateMap = 11'd344;
    356: stateMap = 11'd345;
    357: stateMap = 11'd346;
    358: stateMap = 11'd317;
    359: stateMap = 11'd347;
    360: stateMap = 11'd348;
    361: stateMap = 11'd349;
    362: stateMap = 11'd350;
    363: stateMap = 11'd351;
    364: stateMap = 11'd352;
    365: stateMap = 11'd353;
    366: stateMap = 11'd354;
    367: stateMap = 11'd355;
    368: stateMap = 11'd356;
    369: stateMap = 11'd357;
    370: stateMap = 11'd358;
    371: stateMap = 11'd359;
    372: stateMap = 11'd360;
    373: stateMap = 11'd361;
    374: stateMap = 11'd362;
    375: stateMap = 11'd363;
    376: stateMap = 11'd364;
    377: stateMap = 11'd365;
    378: stateMap = 11'd366;
    379: stateMap = 11'd367;
    380: stateMap = 11'd368;
    381: stateMap = 11'd369;
    382: stateMap = 11'd370;
    383: stateMap = 11'd371;
    384: stateMap = 11'd372;
    385: stateMap = 11'd373;
    386: stateMap = 11'd374;
    387: stateMap = 11'd375;
    388: stateMap = 11'd376;
    389: stateMap = 11'd377;
    390: stateMap = 11'd378;
    391: stateMap = 11'd379;
    392: stateMap = 11'd380;
    393: stateMap = 11'd356;
    394: stateMap = 11'd381;
    395: stateMap = 11'd382;
    396: stateMap = 11'd383;
    397: stateMap = 11'd384;
    398: stateMap = 11'd385;
    399: stateMap = 11'd386;
    400: stateMap = 11'd387;
    401: stateMap = 11'd388;
    402: stateMap = 11'd389;
    403: stateMap = 11'd390;
    404: stateMap = 11'd391;
    405: stateMap = 11'd392;
    406: stateMap = 11'd393;
    407: stateMap = 11'd394;
    408: stateMap = 11'd395;
    409: stateMap = 11'd396;
    410: stateMap = 11'd397;
    411: stateMap = 11'd398;
    412: stateMap = 11'd399;
    413: stateMap = 11'd400;
    414: stateMap = 11'd401;
    415: stateMap = 11'd402;
    416: stateMap = 11'd403;
    417: stateMap = 11'd404;
    418: stateMap = 11'd405;
    419: stateMap = 11'd406;
    420: stateMap = 11'd407;
    421: stateMap = 11'd385;
    422: stateMap = 11'd408;
    423: stateMap = 11'd409;
    424: stateMap = 11'd410;
    425: stateMap = 11'd411;
    426: stateMap = 11'd412;
    427: stateMap = 11'd413;
    428: stateMap = 11'd414;
    429: stateMap = 11'd415;
    430: stateMap = 11'd416;
    431: stateMap = 11'd417;
    432: stateMap = 11'd418;
    433: stateMap = 11'd419;
    434: stateMap = 11'd420;
    435: stateMap = 11'd421;
    436: stateMap = 11'd422;
    437: stateMap = 11'd423;
    438: stateMap = 11'd424;
    439: stateMap = 11'd410;
    440: stateMap = 11'd425;
    441: stateMap = 11'd426;
    442: stateMap = 11'd427;
    443: stateMap = 11'd428;
    444: stateMap = 11'd429;
    445: stateMap = 11'd430;
    446: stateMap = 11'd431;
    447: stateMap = 11'd432;
    448: stateMap = 11'd429;
    449: stateMap = 11'd74;
    450: stateMap = 11'd433;
    451: stateMap = 11'd434;
    452: stateMap = 11'd435;
    453: stateMap = 11'd436;
    454: stateMap = 11'd437;
    455: stateMap = 11'd438;
    456: stateMap = 11'd439;
    457: stateMap = 11'd440;
    458: stateMap = 11'd441;
    459: stateMap = 11'd442;
    460: stateMap = 11'd428;
    461: stateMap = 11'd443;
    462: stateMap = 11'd444;
    463: stateMap = 11'd445;
    464: stateMap = 11'd446;
    465: stateMap = 11'd447;
    466: stateMap = 11'd448;
    467: stateMap = 11'd449;
    468: stateMap = 11'd4;
    469: stateMap = 11'd450;
    470: stateMap = 11'd451;
    471: stateMap = 11'd452;
    472: stateMap = 11'd453;
    473: stateMap = 11'd454;
    474: stateMap = 11'd455;
    475: stateMap = 11'd456;
    476: stateMap = 11'd457;
    477: stateMap = 11'd458;
    478: stateMap = 11'd459;
    479: stateMap = 11'd460;
    480: stateMap = 11'd453;
    481: stateMap = 11'd461;
    482: stateMap = 11'd462;
    483: stateMap = 11'd463;
    484: stateMap = 11'd464;
    485: stateMap = 11'd465;
    486: stateMap = 11'd466;
    487: stateMap = 11'd467;
    488: stateMap = 11'd468;
    489: stateMap = 11'd469;
    490: stateMap = 11'd470;
    491: stateMap = 11'd471;
    492: stateMap = 11'd13;
    493: stateMap = 11'd472;
    494: stateMap = 11'd473;
    495: stateMap = 11'd474;
    496: stateMap = 11'd475;
    497: stateMap = 11'd476;
    498: stateMap = 11'd477;
    499: stateMap = 11'd478;
    500: stateMap = 11'd479;
    501: stateMap = 11'd480;
    502: stateMap = 11'd481;
    503: stateMap = 11'd21;
    504: stateMap = 11'd482;
    505: stateMap = 11'd483;
    506: stateMap = 11'd484;
    507: stateMap = 11'd485;
    508: stateMap = 11'd486;
    509: stateMap = 11'd487;
    510: stateMap = 11'd488;
    511: stateMap = 11'd489;
    512: stateMap = 11'd490;
    513: stateMap = 11'd491;
    514: stateMap = 11'd492;
    515: stateMap = 11'd493;
    516: stateMap = 11'd494;
    517: stateMap = 11'd495;
    518: stateMap = 11'd496;
    519: stateMap = 11'd497;
    520: stateMap = 11'd498;
    521: stateMap = 11'd499;
    522: stateMap = 11'd500;
    523: stateMap = 11'd501;
    524: stateMap = 11'd502;
    525: stateMap = 11'd503;
    526: stateMap = 11'd504;
    527: stateMap = 11'd505;
    528: stateMap = 11'd506;
    529: stateMap = 11'd507;
    530: stateMap = 11'd508;
    531: stateMap = 11'd509;
    532: stateMap = 11'd510;
    533: stateMap = 11'd511;
    534: stateMap = 11'd512;
    535: stateMap = 11'd513;
    536: stateMap = 11'd514;
    537: stateMap = 11'd515;
    538: stateMap = 11'd516;
    539: stateMap = 11'd517;
    540: stateMap = 11'd518;
    541: stateMap = 11'd519;
    542: stateMap = 11'd520;
    543: stateMap = 11'd521;
    544: stateMap = 11'd522;
    545: stateMap = 11'd523;
    546: stateMap = 11'd524;
    547: stateMap = 11'd525;
    548: stateMap = 11'd526;
    549: stateMap = 11'd527;
    550: stateMap = 11'd528;
    551: stateMap = 11'd529;
    552: stateMap = 11'd530;
    553: stateMap = 11'd531;
    554: stateMap = 11'd532;
    555: stateMap = 11'd533;
    556: stateMap = 11'd534;
    557: stateMap = 11'd535;
    558: stateMap = 11'd536;
    559: stateMap = 11'd537;
    560: stateMap = 11'd538;
    561: stateMap = 11'd539;
    562: stateMap = 11'd540;
    563: stateMap = 11'd541;
    564: stateMap = 11'd542;
    565: stateMap = 11'd543;
    566: stateMap = 11'd544;
    567: stateMap = 11'd545;
    568: stateMap = 11'd546;
    569: stateMap = 11'd547;
    570: stateMap = 11'd548;
    571: stateMap = 11'd549;
    572: stateMap = 11'd550;
    573: stateMap = 11'd551;
    574: stateMap = 11'd552;
    575: stateMap = 11'd553;
    576: stateMap = 11'd554;
    577: stateMap = 11'd555;
    578: stateMap = 11'd556;
    579: stateMap = 11'd557;
    580: stateMap = 11'd558;
    581: stateMap = 11'd559;
    582: stateMap = 11'd560;
    583: stateMap = 11'd561;
    584: stateMap = 11'd562;
    585: stateMap = 11'd563;
    586: stateMap = 11'd564;
    587: stateMap = 11'd565;
    588: stateMap = 11'd566;
    589: stateMap = 11'd567;
    590: stateMap = 11'd568;
    591: stateMap = 11'd569;
    592: stateMap = 11'd570;
    593: stateMap = 11'd571;
    594: stateMap = 11'd572;
    595: stateMap = 11'd573;
    596: stateMap = 11'd574;
    597: stateMap = 11'd575;
    598: stateMap = 11'd576;
    599: stateMap = 11'd577;
    600: stateMap = 11'd578;
    601: stateMap = 11'd579;
    602: stateMap = 11'd580;
    603: stateMap = 11'd581;
    604: stateMap = 11'd582;
    605: stateMap = 11'd583;
    606: stateMap = 11'd584;
    607: stateMap = 11'd585;
    608: stateMap = 11'd586;
    609: stateMap = 11'd587;
    610: stateMap = 11'd588;
    611: stateMap = 11'd589;
    612: stateMap = 11'd590;
    613: stateMap = 11'd591;
    614: stateMap = 11'd592;
    615: stateMap = 11'd593;
    616: stateMap = 11'd594;
    617: stateMap = 11'd595;
    618: stateMap = 11'd596;
    619: stateMap = 11'd597;
    620: stateMap = 11'd598;
    621: stateMap = 11'd599;
    622: stateMap = 11'd600;
    623: stateMap = 11'd601;
    624: stateMap = 11'd602;
    625: stateMap = 11'd603;
    626: stateMap = 11'd604;
    627: stateMap = 11'd605;
    628: stateMap = 11'd606;
    629: stateMap = 11'd607;
    630: stateMap = 11'd608;
    631: stateMap = 11'd609;
    632: stateMap = 11'd610;
    633: stateMap = 11'd611;
    634: stateMap = 11'd612;
    635: stateMap = 11'd613;
    636: stateMap = 11'd614;
    637: stateMap = 11'd615;
    638: stateMap = 11'd616;
    639: stateMap = 11'd617;
    640: stateMap = 11'd618;
    641: stateMap = 11'd619;
    642: stateMap = 11'd620;
    643: stateMap = 11'd621;
    644: stateMap = 11'd622;
    645: stateMap = 11'd623;
    646: stateMap = 11'd624;
    647: stateMap = 11'd625;
    648: stateMap = 11'd626;
    649: stateMap = 11'd627;
    650: stateMap = 11'd628;
    651: stateMap = 11'd629;
    652: stateMap = 11'd630;
    653: stateMap = 11'd631;
    654: stateMap = 11'd632;
    655: stateMap = 11'd633;
    656: stateMap = 11'd634;
    657: stateMap = 11'd635;
    658: stateMap = 11'd636;
    659: stateMap = 11'd637;
    660: stateMap = 11'd638;
    661: stateMap = 11'd639;
    662: stateMap = 11'd640;
    663: stateMap = 11'd641;
    664: stateMap = 11'd642;
    665: stateMap = 11'd643;
    666: stateMap = 11'd644;
    667: stateMap = 11'd645;
    668: stateMap = 11'd646;
    669: stateMap = 11'd647;
    670: stateMap = 11'd648;
    671: stateMap = 11'd649;
    672: stateMap = 11'd650;
    673: stateMap = 11'd651;
    674: stateMap = 11'd652;
    675: stateMap = 11'd653;
    676: stateMap = 11'd654;
    677: stateMap = 11'd655;
    678: stateMap = 11'd656;
    679: stateMap = 11'd657;
    680: stateMap = 11'd658;
    681: stateMap = 11'd659;
    682: stateMap = 11'd660;
    683: stateMap = 11'd661;
    684: stateMap = 11'd662;
    685: stateMap = 11'd663;
    686: stateMap = 11'd664;
    687: stateMap = 11'd665;
    688: stateMap = 11'd666;
    689: stateMap = 11'd667;
    690: stateMap = 11'd668;
    691: stateMap = 11'd669;
    692: stateMap = 11'd670;
    693: stateMap = 11'd671;
    694: stateMap = 11'd672;
    695: stateMap = 11'd673;
    696: stateMap = 11'd674;
    697: stateMap = 11'd675;
    698: stateMap = 11'd676;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b1;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b1;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b1;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b1;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b1;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b1;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b1;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b1;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b1;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b1;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b0;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b0;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b1;
    62: acceptStates = 1'b0;
    63: acceptStates = 1'b0;
    64: acceptStates = 1'b0;
    65: acceptStates = 1'b0;
    66: acceptStates = 1'b0;
    67: acceptStates = 1'b1;
    68: acceptStates = 1'b1;
    69: acceptStates = 1'b0;
    70: acceptStates = 1'b0;
    71: acceptStates = 1'b0;
    72: acceptStates = 1'b0;
    73: acceptStates = 1'b0;
    74: acceptStates = 1'b0;
    75: acceptStates = 1'b0;
    76: acceptStates = 1'b0;
    77: acceptStates = 1'b1;
    78: acceptStates = 1'b0;
    79: acceptStates = 1'b0;
    80: acceptStates = 1'b0;
    81: acceptStates = 1'b1;
    82: acceptStates = 1'b0;
    83: acceptStates = 1'b0;
    84: acceptStates = 1'b0;
    85: acceptStates = 1'b0;
    86: acceptStates = 1'b0;
    87: acceptStates = 1'b0;
    88: acceptStates = 1'b0;
    89: acceptStates = 1'b0;
    90: acceptStates = 1'b0;
    91: acceptStates = 1'b0;
    92: acceptStates = 1'b0;
    93: acceptStates = 1'b0;
    94: acceptStates = 1'b0;
    95: acceptStates = 1'b0;
    96: acceptStates = 1'b0;
    97: acceptStates = 1'b0;
    98: acceptStates = 1'b0;
    99: acceptStates = 1'b0;
    100: acceptStates = 1'b0;
    101: acceptStates = 1'b0;
    102: acceptStates = 1'b0;
    103: acceptStates = 1'b0;
    104: acceptStates = 1'b0;
    105: acceptStates = 1'b0;
    106: acceptStates = 1'b0;
    107: acceptStates = 1'b0;
    108: acceptStates = 1'b0;
    109: acceptStates = 1'b0;
    110: acceptStates = 1'b0;
    111: acceptStates = 1'b0;
    112: acceptStates = 1'b0;
    113: acceptStates = 1'b0;
    114: acceptStates = 1'b0;
    115: acceptStates = 1'b0;
    116: acceptStates = 1'b0;
    117: acceptStates = 1'b0;
    118: acceptStates = 1'b0;
    119: acceptStates = 1'b0;
    120: acceptStates = 1'b0;
    121: acceptStates = 1'b0;
    122: acceptStates = 1'b0;
    123: acceptStates = 1'b0;
    124: acceptStates = 1'b0;
    125: acceptStates = 1'b1;
    126: acceptStates = 1'b0;
    127: acceptStates = 1'b1;
    128: acceptStates = 1'b0;
    129: acceptStates = 1'b0;
    130: acceptStates = 1'b1;
    131: acceptStates = 1'b0;
    132: acceptStates = 1'b0;
    133: acceptStates = 1'b0;
    134: acceptStates = 1'b0;
    135: acceptStates = 1'b0;
    136: acceptStates = 1'b0;
    137: acceptStates = 1'b0;
    138: acceptStates = 1'b0;
    139: acceptStates = 1'b0;
    140: acceptStates = 1'b0;
    141: acceptStates = 1'b0;
    142: acceptStates = 1'b0;
    143: acceptStates = 1'b0;
    144: acceptStates = 1'b0;
    145: acceptStates = 1'b0;
    146: acceptStates = 1'b0;
    147: acceptStates = 1'b0;
    148: acceptStates = 1'b0;
    149: acceptStates = 1'b0;
    150: acceptStates = 1'b0;
    151: acceptStates = 1'b0;
    152: acceptStates = 1'b0;
    153: acceptStates = 1'b0;
    154: acceptStates = 1'b0;
    155: acceptStates = 1'b0;
    156: acceptStates = 1'b0;
    157: acceptStates = 1'b0;
    158: acceptStates = 1'b0;
    159: acceptStates = 1'b0;
    160: acceptStates = 1'b0;
    161: acceptStates = 1'b0;
    162: acceptStates = 1'b0;
    163: acceptStates = 1'b0;
    164: acceptStates = 1'b0;
    165: acceptStates = 1'b0;
    166: acceptStates = 1'b0;
    167: acceptStates = 1'b0;
    168: acceptStates = 1'b0;
    169: acceptStates = 1'b1;
    170: acceptStates = 1'b0;
    171: acceptStates = 1'b0;
    172: acceptStates = 1'b0;
    173: acceptStates = 1'b0;
    174: acceptStates = 1'b0;
    175: acceptStates = 1'b0;
    176: acceptStates = 1'b0;
    177: acceptStates = 1'b0;
    178: acceptStates = 1'b0;
    179: acceptStates = 1'b0;
    180: acceptStates = 1'b0;
    181: acceptStates = 1'b0;
    182: acceptStates = 1'b0;
    183: acceptStates = 1'b0;
    184: acceptStates = 1'b0;
    185: acceptStates = 1'b0;
    186: acceptStates = 1'b0;
    187: acceptStates = 1'b0;
    188: acceptStates = 1'b0;
    189: acceptStates = 1'b0;
    190: acceptStates = 1'b0;
    191: acceptStates = 1'b0;
    192: acceptStates = 1'b0;
    193: acceptStates = 1'b0;
    194: acceptStates = 1'b0;
    195: acceptStates = 1'b0;
    196: acceptStates = 1'b0;
    197: acceptStates = 1'b0;
    198: acceptStates = 1'b0;
    199: acceptStates = 1'b0;
    200: acceptStates = 1'b0;
    201: acceptStates = 1'b0;
    202: acceptStates = 1'b0;
    203: acceptStates = 1'b0;
    204: acceptStates = 1'b0;
    205: acceptStates = 1'b0;
    206: acceptStates = 1'b1;
    207: acceptStates = 1'b0;
    208: acceptStates = 1'b0;
    209: acceptStates = 1'b0;
    210: acceptStates = 1'b0;
    211: acceptStates = 1'b0;
    212: acceptStates = 1'b0;
    213: acceptStates = 1'b0;
    214: acceptStates = 1'b0;
    215: acceptStates = 1'b0;
    216: acceptStates = 1'b0;
    217: acceptStates = 1'b0;
    218: acceptStates = 1'b0;
    219: acceptStates = 1'b0;
    220: acceptStates = 1'b0;
    221: acceptStates = 1'b0;
    222: acceptStates = 1'b0;
    223: acceptStates = 1'b0;
    224: acceptStates = 1'b0;
    225: acceptStates = 1'b0;
    226: acceptStates = 1'b0;
    227: acceptStates = 1'b0;
    228: acceptStates = 1'b0;
    229: acceptStates = 1'b0;
    230: acceptStates = 1'b0;
    231: acceptStates = 1'b0;
    232: acceptStates = 1'b0;
    233: acceptStates = 1'b0;
    234: acceptStates = 1'b0;
    235: acceptStates = 1'b0;
    236: acceptStates = 1'b0;
    237: acceptStates = 1'b0;
    238: acceptStates = 1'b0;
    239: acceptStates = 1'b0;
    240: acceptStates = 1'b0;
    241: acceptStates = 1'b0;
    242: acceptStates = 1'b0;
    243: acceptStates = 1'b0;
    244: acceptStates = 1'b0;
    245: acceptStates = 1'b0;
    246: acceptStates = 1'b0;
    247: acceptStates = 1'b0;
    248: acceptStates = 1'b0;
    249: acceptStates = 1'b0;
    250: acceptStates = 1'b0;
    251: acceptStates = 1'b1;
    252: acceptStates = 1'b0;
    253: acceptStates = 1'b0;
    254: acceptStates = 1'b0;
    255: acceptStates = 1'b0;
    256: acceptStates = 1'b0;
    257: acceptStates = 1'b0;
    258: acceptStates = 1'b0;
    259: acceptStates = 1'b0;
    260: acceptStates = 1'b0;
    261: acceptStates = 1'b0;
    262: acceptStates = 1'b0;
    263: acceptStates = 1'b0;
    264: acceptStates = 1'b0;
    265: acceptStates = 1'b0;
    266: acceptStates = 1'b0;
    267: acceptStates = 1'b0;
    268: acceptStates = 1'b0;
    269: acceptStates = 1'b0;
    270: acceptStates = 1'b0;
    271: acceptStates = 1'b0;
    272: acceptStates = 1'b0;
    273: acceptStates = 1'b0;
    274: acceptStates = 1'b0;
    275: acceptStates = 1'b0;
    276: acceptStates = 1'b0;
    277: acceptStates = 1'b0;
    278: acceptStates = 1'b0;
    279: acceptStates = 1'b0;
    280: acceptStates = 1'b0;
    281: acceptStates = 1'b0;
    282: acceptStates = 1'b0;
    283: acceptStates = 1'b0;
    284: acceptStates = 1'b0;
    285: acceptStates = 1'b0;
    286: acceptStates = 1'b0;
    287: acceptStates = 1'b0;
    288: acceptStates = 1'b0;
    289: acceptStates = 1'b0;
    290: acceptStates = 1'b0;
    291: acceptStates = 1'b1;
    292: acceptStates = 1'b0;
    293: acceptStates = 1'b0;
    294: acceptStates = 1'b0;
    295: acceptStates = 1'b0;
    296: acceptStates = 1'b0;
    297: acceptStates = 1'b0;
    298: acceptStates = 1'b0;
    299: acceptStates = 1'b0;
    300: acceptStates = 1'b0;
    301: acceptStates = 1'b0;
    302: acceptStates = 1'b0;
    303: acceptStates = 1'b0;
    304: acceptStates = 1'b0;
    305: acceptStates = 1'b0;
    306: acceptStates = 1'b0;
    307: acceptStates = 1'b0;
    308: acceptStates = 1'b0;
    309: acceptStates = 1'b0;
    310: acceptStates = 1'b0;
    311: acceptStates = 1'b0;
    312: acceptStates = 1'b0;
    313: acceptStates = 1'b0;
    314: acceptStates = 1'b0;
    315: acceptStates = 1'b0;
    316: acceptStates = 1'b0;
    317: acceptStates = 1'b0;
    318: acceptStates = 1'b0;
    319: acceptStates = 1'b0;
    320: acceptStates = 1'b0;
    321: acceptStates = 1'b0;
    322: acceptStates = 1'b0;
    323: acceptStates = 1'b0;
    324: acceptStates = 1'b0;
    325: acceptStates = 1'b0;
    326: acceptStates = 1'b0;
    327: acceptStates = 1'b0;
    328: acceptStates = 1'b1;
    329: acceptStates = 1'b0;
    330: acceptStates = 1'b0;
    331: acceptStates = 1'b0;
    332: acceptStates = 1'b0;
    333: acceptStates = 1'b0;
    334: acceptStates = 1'b0;
    335: acceptStates = 1'b0;
    336: acceptStates = 1'b0;
    337: acceptStates = 1'b0;
    338: acceptStates = 1'b0;
    339: acceptStates = 1'b0;
    340: acceptStates = 1'b0;
    341: acceptStates = 1'b0;
    342: acceptStates = 1'b0;
    343: acceptStates = 1'b0;
    344: acceptStates = 1'b0;
    345: acceptStates = 1'b0;
    346: acceptStates = 1'b0;
    347: acceptStates = 1'b0;
    348: acceptStates = 1'b0;
    349: acceptStates = 1'b0;
    350: acceptStates = 1'b0;
    351: acceptStates = 1'b0;
    352: acceptStates = 1'b0;
    353: acceptStates = 1'b0;
    354: acceptStates = 1'b0;
    355: acceptStates = 1'b0;
    356: acceptStates = 1'b0;
    357: acceptStates = 1'b0;
    358: acceptStates = 1'b0;
    359: acceptStates = 1'b0;
    360: acceptStates = 1'b0;
    361: acceptStates = 1'b0;
    362: acceptStates = 1'b0;
    363: acceptStates = 1'b0;
    364: acceptStates = 1'b0;
    365: acceptStates = 1'b0;
    366: acceptStates = 1'b0;
    367: acceptStates = 1'b0;
    368: acceptStates = 1'b1;
    369: acceptStates = 1'b0;
    370: acceptStates = 1'b0;
    371: acceptStates = 1'b0;
    372: acceptStates = 1'b0;
    373: acceptStates = 1'b0;
    374: acceptStates = 1'b0;
    375: acceptStates = 1'b0;
    376: acceptStates = 1'b0;
    377: acceptStates = 1'b0;
    378: acceptStates = 1'b0;
    379: acceptStates = 1'b0;
    380: acceptStates = 1'b0;
    381: acceptStates = 1'b0;
    382: acceptStates = 1'b0;
    383: acceptStates = 1'b0;
    384: acceptStates = 1'b0;
    385: acceptStates = 1'b0;
    386: acceptStates = 1'b0;
    387: acceptStates = 1'b0;
    388: acceptStates = 1'b0;
    389: acceptStates = 1'b0;
    390: acceptStates = 1'b0;
    391: acceptStates = 1'b0;
    392: acceptStates = 1'b0;
    393: acceptStates = 1'b0;
    394: acceptStates = 1'b0;
    395: acceptStates = 1'b0;
    396: acceptStates = 1'b0;
    397: acceptStates = 1'b0;
    398: acceptStates = 1'b1;
    399: acceptStates = 1'b0;
    400: acceptStates = 1'b0;
    401: acceptStates = 1'b0;
    402: acceptStates = 1'b0;
    403: acceptStates = 1'b0;
    404: acceptStates = 1'b0;
    405: acceptStates = 1'b0;
    406: acceptStates = 1'b0;
    407: acceptStates = 1'b0;
    408: acceptStates = 1'b0;
    409: acceptStates = 1'b0;
    410: acceptStates = 1'b0;
    411: acceptStates = 1'b0;
    412: acceptStates = 1'b0;
    413: acceptStates = 1'b0;
    414: acceptStates = 1'b0;
    415: acceptStates = 1'b0;
    416: acceptStates = 1'b0;
    417: acceptStates = 1'b0;
    418: acceptStates = 1'b0;
    419: acceptStates = 1'b0;
    420: acceptStates = 1'b0;
    421: acceptStates = 1'b0;
    422: acceptStates = 1'b0;
    423: acceptStates = 1'b0;
    424: acceptStates = 1'b1;
    425: acceptStates = 1'b0;
    426: acceptStates = 1'b0;
    427: acceptStates = 1'b0;
    428: acceptStates = 1'b0;
    429: acceptStates = 1'b0;
    430: acceptStates = 1'b0;
    431: acceptStates = 1'b0;
    432: acceptStates = 1'b0;
    433: acceptStates = 1'b0;
    434: acceptStates = 1'b0;
    435: acceptStates = 1'b0;
    436: acceptStates = 1'b0;
    437: acceptStates = 1'b0;
    438: acceptStates = 1'b0;
    439: acceptStates = 1'b0;
    440: acceptStates = 1'b0;
    441: acceptStates = 1'b0;
    442: acceptStates = 1'b0;
    443: acceptStates = 1'b1;
    444: acceptStates = 1'b0;
    445: acceptStates = 1'b0;
    446: acceptStates = 1'b0;
    447: acceptStates = 1'b0;
    448: acceptStates = 1'b1;
    449: acceptStates = 1'b0;
    450: acceptStates = 1'b0;
    451: acceptStates = 1'b0;
    452: acceptStates = 1'b0;
    453: acceptStates = 1'b0;
    454: acceptStates = 1'b0;
    455: acceptStates = 1'b0;
    456: acceptStates = 1'b0;
    457: acceptStates = 1'b0;
    458: acceptStates = 1'b0;
    459: acceptStates = 1'b0;
    460: acceptStates = 1'b0;
    461: acceptStates = 1'b0;
    462: acceptStates = 1'b0;
    463: acceptStates = 1'b0;
    464: acceptStates = 1'b0;
    465: acceptStates = 1'b0;
    466: acceptStates = 1'b0;
    467: acceptStates = 1'b0;
    468: acceptStates = 1'b0;
    469: acceptStates = 1'b0;
    470: acceptStates = 1'b0;
    471: acceptStates = 1'b0;
    472: acceptStates = 1'b1;
    473: acceptStates = 1'b0;
    474: acceptStates = 1'b0;
    475: acceptStates = 1'b0;
    476: acceptStates = 1'b0;
    477: acceptStates = 1'b0;
    478: acceptStates = 1'b0;
    479: acceptStates = 1'b0;
    480: acceptStates = 1'b0;
    481: acceptStates = 1'b0;
    482: acceptStates = 1'b0;
    483: acceptStates = 1'b0;
    484: acceptStates = 1'b0;
    485: acceptStates = 1'b0;
    486: acceptStates = 1'b0;
    487: acceptStates = 1'b0;
    488: acceptStates = 1'b0;
    489: acceptStates = 1'b0;
    490: acceptStates = 1'b0;
    491: acceptStates = 1'b0;
    492: acceptStates = 1'b1;
    493: acceptStates = 1'b0;
    494: acceptStates = 1'b0;
    495: acceptStates = 1'b0;
    496: acceptStates = 1'b0;
    497: acceptStates = 1'b0;
    498: acceptStates = 1'b0;
    499: acceptStates = 1'b0;
    500: acceptStates = 1'b0;
    501: acceptStates = 1'b0;
    502: acceptStates = 1'b0;
    503: acceptStates = 1'b0;
    504: acceptStates = 1'b0;
    505: acceptStates = 1'b0;
    506: acceptStates = 1'b0;
    507: acceptStates = 1'b0;
    508: acceptStates = 1'b0;
    509: acceptStates = 1'b0;
    510: acceptStates = 1'b0;
    511: acceptStates = 1'b0;
    512: acceptStates = 1'b0;
    513: acceptStates = 1'b0;
    514: acceptStates = 1'b0;
    515: acceptStates = 1'b0;
    516: acceptStates = 1'b0;
    517: acceptStates = 1'b0;
    518: acceptStates = 1'b0;
    519: acceptStates = 1'b0;
    520: acceptStates = 1'b0;
    521: acceptStates = 1'b0;
    522: acceptStates = 1'b0;
    523: acceptStates = 1'b0;
    524: acceptStates = 1'b0;
    525: acceptStates = 1'b0;
    526: acceptStates = 1'b0;
    527: acceptStates = 1'b0;
    528: acceptStates = 1'b0;
    529: acceptStates = 1'b0;
    530: acceptStates = 1'b0;
    531: acceptStates = 1'b0;
    532: acceptStates = 1'b0;
    533: acceptStates = 1'b0;
    534: acceptStates = 1'b0;
    535: acceptStates = 1'b0;
    536: acceptStates = 1'b0;
    537: acceptStates = 1'b0;
    538: acceptStates = 1'b0;
    539: acceptStates = 1'b0;
    540: acceptStates = 1'b0;
    541: acceptStates = 1'b0;
    542: acceptStates = 1'b0;
    543: acceptStates = 1'b0;
    544: acceptStates = 1'b0;
    545: acceptStates = 1'b0;
    546: acceptStates = 1'b0;
    547: acceptStates = 1'b0;
    548: acceptStates = 1'b0;
    549: acceptStates = 1'b0;
    550: acceptStates = 1'b0;
    551: acceptStates = 1'b0;
    552: acceptStates = 1'b0;
    553: acceptStates = 1'b0;
    554: acceptStates = 1'b0;
    555: acceptStates = 1'b0;
    556: acceptStates = 1'b0;
    557: acceptStates = 1'b0;
    558: acceptStates = 1'b0;
    559: acceptStates = 1'b0;
    560: acceptStates = 1'b0;
    561: acceptStates = 1'b0;
    562: acceptStates = 1'b0;
    563: acceptStates = 1'b0;
    564: acceptStates = 1'b0;
    565: acceptStates = 1'b0;
    566: acceptStates = 1'b0;
    567: acceptStates = 1'b0;
    568: acceptStates = 1'b0;
    569: acceptStates = 1'b0;
    570: acceptStates = 1'b0;
    571: acceptStates = 1'b0;
    572: acceptStates = 1'b0;
    573: acceptStates = 1'b0;
    574: acceptStates = 1'b0;
    575: acceptStates = 1'b0;
    576: acceptStates = 1'b0;
    577: acceptStates = 1'b0;
    578: acceptStates = 1'b0;
    579: acceptStates = 1'b0;
    580: acceptStates = 1'b0;
    581: acceptStates = 1'b0;
    582: acceptStates = 1'b0;
    583: acceptStates = 1'b0;
    584: acceptStates = 1'b0;
    585: acceptStates = 1'b0;
    586: acceptStates = 1'b0;
    587: acceptStates = 1'b0;
    588: acceptStates = 1'b0;
    589: acceptStates = 1'b0;
    590: acceptStates = 1'b0;
    591: acceptStates = 1'b0;
    592: acceptStates = 1'b0;
    593: acceptStates = 1'b0;
    594: acceptStates = 1'b0;
    595: acceptStates = 1'b0;
    596: acceptStates = 1'b0;
    597: acceptStates = 1'b0;
    598: acceptStates = 1'b0;
    599: acceptStates = 1'b0;
    600: acceptStates = 1'b0;
    601: acceptStates = 1'b0;
    602: acceptStates = 1'b0;
    603: acceptStates = 1'b0;
    604: acceptStates = 1'b0;
    605: acceptStates = 1'b0;
    606: acceptStates = 1'b0;
    607: acceptStates = 1'b0;
    608: acceptStates = 1'b0;
    609: acceptStates = 1'b0;
    610: acceptStates = 1'b0;
    611: acceptStates = 1'b0;
    612: acceptStates = 1'b0;
    613: acceptStates = 1'b0;
    614: acceptStates = 1'b0;
    615: acceptStates = 1'b0;
    616: acceptStates = 1'b0;
    617: acceptStates = 1'b0;
    618: acceptStates = 1'b0;
    619: acceptStates = 1'b0;
    620: acceptStates = 1'b0;
    621: acceptStates = 1'b0;
    622: acceptStates = 1'b0;
    623: acceptStates = 1'b0;
    624: acceptStates = 1'b0;
    625: acceptStates = 1'b0;
    626: acceptStates = 1'b0;
    627: acceptStates = 1'b0;
    628: acceptStates = 1'b0;
    629: acceptStates = 1'b0;
    630: acceptStates = 1'b0;
    631: acceptStates = 1'b0;
    632: acceptStates = 1'b0;
    633: acceptStates = 1'b0;
    634: acceptStates = 1'b0;
    635: acceptStates = 1'b0;
    636: acceptStates = 1'b0;
    637: acceptStates = 1'b0;
    638: acceptStates = 1'b0;
    639: acceptStates = 1'b0;
    640: acceptStates = 1'b0;
    641: acceptStates = 1'b0;
    642: acceptStates = 1'b0;
    643: acceptStates = 1'b0;
    644: acceptStates = 1'b0;
    645: acceptStates = 1'b0;
    646: acceptStates = 1'b0;
    647: acceptStates = 1'b0;
    648: acceptStates = 1'b0;
    649: acceptStates = 1'b0;
    650: acceptStates = 1'b0;
    651: acceptStates = 1'b0;
    652: acceptStates = 1'b0;
    653: acceptStates = 1'b0;
    654: acceptStates = 1'b0;
    655: acceptStates = 1'b0;
    656: acceptStates = 1'b0;
    657: acceptStates = 1'b0;
    658: acceptStates = 1'b0;
    659: acceptStates = 1'b0;
    660: acceptStates = 1'b0;
    661: acceptStates = 1'b0;
    662: acceptStates = 1'b0;
    663: acceptStates = 1'b0;
    664: acceptStates = 1'b0;
    665: acceptStates = 1'b0;
    666: acceptStates = 1'b0;
    667: acceptStates = 1'b0;
    668: acceptStates = 1'b0;
    669: acceptStates = 1'b0;
    670: acceptStates = 1'b0;
    671: acceptStates = 1'b0;
    672: acceptStates = 1'b0;
    673: acceptStates = 1'b0;
    674: acceptStates = 1'b0;
    675: acceptStates = 1'b0;
    676: acceptStates = 1'b0;
    677: acceptStates = 1'b0;
    678: acceptStates = 1'b0;
    679: acceptStates = 1'b0;
    680: acceptStates = 1'b0;
    681: acceptStates = 1'b0;
    682: acceptStates = 1'b0;
    683: acceptStates = 1'b0;
    684: acceptStates = 1'b0;
    685: acceptStates = 1'b0;
    686: acceptStates = 1'b0;
    687: acceptStates = 1'b0;
    688: acceptStates = 1'b0;
    689: acceptStates = 1'b0;
    690: acceptStates = 1'b0;
    691: acceptStates = 1'b0;
    692: acceptStates = 1'b0;
    693: acceptStates = 1'b0;
    694: acceptStates = 1'b0;
    695: acceptStates = 1'b0;
    696: acceptStates = 1'b0;
    697: acceptStates = 1'b0;
    698: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd1;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd124;
      3: stateTransition = 11'd124;
      4: stateTransition = 11'd124;
      5: stateTransition = 11'd124;
      6: stateTransition = 11'd124;
      7: stateTransition = 11'd124;
      8: stateTransition = 11'd124;
      9: stateTransition = 11'd124;
      10: stateTransition = 11'd124;
      11: stateTransition = 11'd124;
      12: stateTransition = 11'd124;
      13: stateTransition = 11'd124;
      14: stateTransition = 11'd124;
      15: stateTransition = 11'd124;
      16: stateTransition = 11'd124;
      17: stateTransition = 11'd124;
      18: stateTransition = 11'd124;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd124;
      22: stateTransition = 11'd124;
      23: stateTransition = 11'd124;
      24: stateTransition = 11'd124;
      25: stateTransition = 11'd124;
      26: stateTransition = 11'd124;
      27: stateTransition = 11'd124;
      28: stateTransition = 11'd124;
      29: stateTransition = 11'd124;
      30: stateTransition = 11'd124;
      31: stateTransition = 11'd124;
      32: stateTransition = 11'd124;
      33: stateTransition = 11'd124;
      34: stateTransition = 11'd124;
      35: stateTransition = 11'd124;
      36: stateTransition = 11'd124;
      37: stateTransition = 11'd124;
      38: stateTransition = 11'd124;
      39: stateTransition = 11'd124;
      40: stateTransition = 11'd136;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd449;
      2: stateTransition = 11'd449;
      3: stateTransition = 11'd449;
      4: stateTransition = 11'd449;
      5: stateTransition = 11'd449;
      6: stateTransition = 11'd77;
      7: stateTransition = 11'd449;
      8: stateTransition = 11'd449;
      9: stateTransition = 11'd449;
      10: stateTransition = 11'd449;
      11: stateTransition = 11'd449;
      12: stateTransition = 11'd449;
      13: stateTransition = 11'd449;
      14: stateTransition = 11'd449;
      15: stateTransition = 11'd449;
      16: stateTransition = 11'd449;
      17: stateTransition = 11'd449;
      18: stateTransition = 11'd449;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd449;
      22: stateTransition = 11'd449;
      23: stateTransition = 11'd449;
      24: stateTransition = 11'd449;
      25: stateTransition = 11'd449;
      26: stateTransition = 11'd449;
      27: stateTransition = 11'd449;
      28: stateTransition = 11'd449;
      29: stateTransition = 11'd449;
      30: stateTransition = 11'd449;
      31: stateTransition = 11'd449;
      32: stateTransition = 11'd449;
      33: stateTransition = 11'd449;
      34: stateTransition = 11'd449;
      35: stateTransition = 11'd449;
      36: stateTransition = 11'd449;
      37: stateTransition = 11'd449;
      38: stateTransition = 11'd449;
      39: stateTransition = 11'd449;
      40: stateTransition = 11'd449;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd140;
      2: stateTransition = 11'd62;
      3: stateTransition = 11'd140;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd140;
      6: stateTransition = 11'd140;
      7: stateTransition = 11'd140;
      8: stateTransition = 11'd140;
      9: stateTransition = 11'd78;
      10: stateTransition = 11'd140;
      11: stateTransition = 11'd140;
      12: stateTransition = 11'd140;
      13: stateTransition = 11'd140;
      14: stateTransition = 11'd140;
      15: stateTransition = 11'd140;
      16: stateTransition = 11'd140;
      17: stateTransition = 11'd140;
      18: stateTransition = 11'd140;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd140;
      22: stateTransition = 11'd173;
      23: stateTransition = 11'd140;
      24: stateTransition = 11'd140;
      25: stateTransition = 11'd140;
      26: stateTransition = 11'd140;
      27: stateTransition = 11'd140;
      28: stateTransition = 11'd140;
      29: stateTransition = 11'd140;
      30: stateTransition = 11'd140;
      31: stateTransition = 11'd140;
      32: stateTransition = 11'd140;
      33: stateTransition = 11'd140;
      34: stateTransition = 11'd140;
      35: stateTransition = 11'd140;
      36: stateTransition = 11'd140;
      37: stateTransition = 11'd140;
      38: stateTransition = 11'd140;
      39: stateTransition = 11'd140;
      40: stateTransition = 11'd140;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd460;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd460;
      10: stateTransition = 11'd460;
      11: stateTransition = 11'd460;
      12: stateTransition = 11'd460;
      13: stateTransition = 11'd460;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd460;
      16: stateTransition = 11'd460;
      17: stateTransition = 11'd460;
      18: stateTransition = 11'd460;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd460;
      22: stateTransition = 11'd460;
      23: stateTransition = 11'd460;
      24: stateTransition = 11'd460;
      25: stateTransition = 11'd460;
      26: stateTransition = 11'd460;
      27: stateTransition = 11'd460;
      28: stateTransition = 11'd460;
      29: stateTransition = 11'd460;
      30: stateTransition = 11'd460;
      31: stateTransition = 11'd460;
      32: stateTransition = 11'd460;
      33: stateTransition = 11'd460;
      34: stateTransition = 11'd460;
      35: stateTransition = 11'd460;
      36: stateTransition = 11'd460;
      37: stateTransition = 11'd460;
      38: stateTransition = 11'd460;
      39: stateTransition = 11'd460;
      40: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd63;
      2: stateTransition = 11'd63;
      3: stateTransition = 11'd63;
      4: stateTransition = 11'd79;
      5: stateTransition = 11'd63;
      6: stateTransition = 11'd2;
      7: stateTransition = 11'd63;
      8: stateTransition = 11'd63;
      9: stateTransition = 11'd63;
      10: stateTransition = 11'd63;
      11: stateTransition = 11'd63;
      12: stateTransition = 11'd63;
      13: stateTransition = 11'd63;
      14: stateTransition = 11'd63;
      15: stateTransition = 11'd63;
      16: stateTransition = 11'd63;
      17: stateTransition = 11'd63;
      18: stateTransition = 11'd63;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd63;
      22: stateTransition = 11'd63;
      23: stateTransition = 11'd63;
      24: stateTransition = 11'd63;
      25: stateTransition = 11'd63;
      26: stateTransition = 11'd63;
      27: stateTransition = 11'd63;
      28: stateTransition = 11'd63;
      29: stateTransition = 11'd63;
      30: stateTransition = 11'd63;
      31: stateTransition = 11'd63;
      32: stateTransition = 11'd63;
      33: stateTransition = 11'd63;
      34: stateTransition = 11'd63;
      35: stateTransition = 11'd63;
      36: stateTransition = 11'd63;
      37: stateTransition = 11'd63;
      38: stateTransition = 11'd63;
      39: stateTransition = 11'd63;
      40: stateTransition = 11'd63;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd127;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd127;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd127;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd127;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd468;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd4;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd468;
      10: stateTransition = 11'd468;
      11: stateTransition = 11'd468;
      12: stateTransition = 11'd468;
      13: stateTransition = 11'd468;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd468;
      16: stateTransition = 11'd468;
      17: stateTransition = 11'd468;
      18: stateTransition = 11'd468;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd468;
      22: stateTransition = 11'd468;
      23: stateTransition = 11'd468;
      24: stateTransition = 11'd468;
      25: stateTransition = 11'd468;
      26: stateTransition = 11'd468;
      27: stateTransition = 11'd468;
      28: stateTransition = 11'd468;
      29: stateTransition = 11'd468;
      30: stateTransition = 11'd468;
      31: stateTransition = 11'd468;
      32: stateTransition = 11'd468;
      33: stateTransition = 11'd468;
      34: stateTransition = 11'd468;
      35: stateTransition = 11'd468;
      36: stateTransition = 11'd468;
      37: stateTransition = 11'd468;
      38: stateTransition = 11'd468;
      39: stateTransition = 11'd468;
      40: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd27;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd27;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd27;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd445;
      2: stateTransition = 11'd445;
      3: stateTransition = 11'd445;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd456;
      8: stateTransition = 11'd445;
      9: stateTransition = 11'd445;
      10: stateTransition = 11'd445;
      11: stateTransition = 11'd445;
      12: stateTransition = 11'd445;
      13: stateTransition = 11'd654;
      14: stateTransition = 11'd445;
      15: stateTransition = 11'd445;
      16: stateTransition = 11'd445;
      17: stateTransition = 11'd445;
      18: stateTransition = 11'd445;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd445;
      22: stateTransition = 11'd445;
      23: stateTransition = 11'd445;
      24: stateTransition = 11'd445;
      25: stateTransition = 11'd445;
      26: stateTransition = 11'd445;
      27: stateTransition = 11'd445;
      28: stateTransition = 11'd445;
      29: stateTransition = 11'd445;
      30: stateTransition = 11'd445;
      31: stateTransition = 11'd445;
      32: stateTransition = 11'd445;
      33: stateTransition = 11'd445;
      34: stateTransition = 11'd445;
      35: stateTransition = 11'd445;
      36: stateTransition = 11'd445;
      37: stateTransition = 11'd445;
      38: stateTransition = 11'd445;
      39: stateTransition = 11'd445;
      40: stateTransition = 11'd445;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd67;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd67;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd67;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd67;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd426;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd426;
      10: stateTransition = 11'd468;
      11: stateTransition = 11'd426;
      12: stateTransition = 11'd468;
      13: stateTransition = 11'd426;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd4;
      16: stateTransition = 11'd426;
      17: stateTransition = 11'd468;
      18: stateTransition = 11'd426;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd468;
      22: stateTransition = 11'd468;
      23: stateTransition = 11'd468;
      24: stateTransition = 11'd468;
      25: stateTransition = 11'd426;
      26: stateTransition = 11'd468;
      27: stateTransition = 11'd468;
      28: stateTransition = 11'd468;
      29: stateTransition = 11'd426;
      30: stateTransition = 11'd468;
      31: stateTransition = 11'd468;
      32: stateTransition = 11'd426;
      33: stateTransition = 11'd468;
      34: stateTransition = 11'd468;
      35: stateTransition = 11'd468;
      36: stateTransition = 11'd468;
      37: stateTransition = 11'd468;
      38: stateTransition = 11'd468;
      39: stateTransition = 11'd426;
      40: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd17;
      2: stateTransition = 11'd17;
      3: stateTransition = 11'd17;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd17;
      8: stateTransition = 11'd17;
      9: stateTransition = 11'd17;
      10: stateTransition = 11'd17;
      11: stateTransition = 11'd17;
      12: stateTransition = 11'd372;
      13: stateTransition = 11'd539;
      14: stateTransition = 11'd17;
      15: stateTransition = 11'd17;
      16: stateTransition = 11'd17;
      17: stateTransition = 11'd17;
      18: stateTransition = 11'd17;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd17;
      22: stateTransition = 11'd17;
      23: stateTransition = 11'd17;
      24: stateTransition = 11'd17;
      25: stateTransition = 11'd17;
      26: stateTransition = 11'd17;
      27: stateTransition = 11'd17;
      28: stateTransition = 11'd17;
      29: stateTransition = 11'd17;
      30: stateTransition = 11'd17;
      31: stateTransition = 11'd17;
      32: stateTransition = 11'd17;
      33: stateTransition = 11'd17;
      34: stateTransition = 11'd17;
      35: stateTransition = 11'd17;
      36: stateTransition = 11'd17;
      37: stateTransition = 11'd17;
      38: stateTransition = 11'd17;
      39: stateTransition = 11'd17;
      40: stateTransition = 11'd17;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd329;
      2: stateTransition = 11'd329;
      3: stateTransition = 11'd329;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd329;
      8: stateTransition = 11'd329;
      9: stateTransition = 11'd329;
      10: stateTransition = 11'd329;
      11: stateTransition = 11'd329;
      12: stateTransition = 11'd329;
      13: stateTransition = 11'd548;
      14: stateTransition = 11'd329;
      15: stateTransition = 11'd329;
      16: stateTransition = 11'd329;
      17: stateTransition = 11'd329;
      18: stateTransition = 11'd329;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd329;
      22: stateTransition = 11'd329;
      23: stateTransition = 11'd329;
      24: stateTransition = 11'd329;
      25: stateTransition = 11'd329;
      26: stateTransition = 11'd329;
      27: stateTransition = 11'd329;
      28: stateTransition = 11'd329;
      29: stateTransition = 11'd329;
      30: stateTransition = 11'd329;
      31: stateTransition = 11'd329;
      32: stateTransition = 11'd329;
      33: stateTransition = 11'd329;
      34: stateTransition = 11'd329;
      35: stateTransition = 11'd329;
      36: stateTransition = 11'd329;
      37: stateTransition = 11'd329;
      38: stateTransition = 11'd329;
      39: stateTransition = 11'd329;
      40: stateTransition = 11'd329;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd68;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd68;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd68;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd68;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd6;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd6;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd6;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd16;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd16;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd16;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd16;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd25;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd25;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd25;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd25;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd8;
      16: stateTransition = 11'd25;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd25;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd25;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd25;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd25;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd25;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd10;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd10;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd10;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd29;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd29;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd29;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd29;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd12;
      16: stateTransition = 11'd29;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd29;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd29;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd29;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd29;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd29;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd14;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd14;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd14;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd37;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd37;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd37;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd38;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd37;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd38;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd38;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd38;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd38;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd16;
      16: stateTransition = 11'd38;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd38;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd38;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd38;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd38;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd38;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd39;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd39;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd39;
      12: stateTransition = 11'd40;
      13: stateTransition = 11'd39;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd39;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd39;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd39;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd39;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd39;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd39;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd41;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd41;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd41;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd18;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd18;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd18;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd51;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd53;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd37;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd37;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd37;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd38;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd37;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd38;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd38;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd38;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd38;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd16;
      16: stateTransition = 11'd38;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd38;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd38;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd38;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd38;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd38;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd39;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd39;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd39;
      12: stateTransition = 11'd40;
      13: stateTransition = 11'd39;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd39;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd39;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd39;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd39;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd39;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd39;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd41;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd41;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd41;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd73;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd73;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd73;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd73;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd44;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd44;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd44;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd74;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd74;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd74;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd74;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd47;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd47;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd47;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd75;
      17: stateTransition = 11'd48;
      18: stateTransition = 11'd75;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd75;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd75;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd48;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd76;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd76;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd76;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd51;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd76;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd18;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd18;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd18;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd51;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd54;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd16;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd22;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd22;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd492;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd472;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd492;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd492;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd181;
      2: stateTransition = 11'd181;
      3: stateTransition = 11'd5;
      4: stateTransition = 11'd181;
      5: stateTransition = 11'd181;
      6: stateTransition = 11'd181;
      7: stateTransition = 11'd217;
      8: stateTransition = 11'd181;
      9: stateTransition = 11'd181;
      10: stateTransition = 11'd181;
      11: stateTransition = 11'd181;
      12: stateTransition = 11'd181;
      13: stateTransition = 11'd181;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd181;
      16: stateTransition = 11'd181;
      17: stateTransition = 11'd181;
      18: stateTransition = 11'd181;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd181;
      22: stateTransition = 11'd181;
      23: stateTransition = 11'd181;
      24: stateTransition = 11'd181;
      25: stateTransition = 11'd181;
      26: stateTransition = 11'd181;
      27: stateTransition = 11'd181;
      28: stateTransition = 11'd181;
      29: stateTransition = 11'd181;
      30: stateTransition = 11'd181;
      31: stateTransition = 11'd181;
      32: stateTransition = 11'd181;
      33: stateTransition = 11'd181;
      34: stateTransition = 11'd181;
      35: stateTransition = 11'd181;
      36: stateTransition = 11'd181;
      37: stateTransition = 11'd181;
      38: stateTransition = 11'd181;
      39: stateTransition = 11'd181;
      40: stateTransition = 11'd181;
      default: stateTransition = 11'bX;
    endcase
    60: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd7;
      2: stateTransition = 11'd7;
      3: stateTransition = 11'd7;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd7;
      6: stateTransition = 11'd61;
      7: stateTransition = 11'd7;
      8: stateTransition = 11'd7;
      9: stateTransition = 11'd7;
      10: stateTransition = 11'd7;
      11: stateTransition = 11'd7;
      12: stateTransition = 11'd7;
      13: stateTransition = 11'd7;
      14: stateTransition = 11'd7;
      15: stateTransition = 11'd7;
      16: stateTransition = 11'd7;
      17: stateTransition = 11'd7;
      18: stateTransition = 11'd7;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd7;
      22: stateTransition = 11'd7;
      23: stateTransition = 11'd7;
      24: stateTransition = 11'd7;
      25: stateTransition = 11'd7;
      26: stateTransition = 11'd7;
      27: stateTransition = 11'd7;
      28: stateTransition = 11'd7;
      29: stateTransition = 11'd7;
      30: stateTransition = 11'd7;
      31: stateTransition = 11'd7;
      32: stateTransition = 11'd7;
      33: stateTransition = 11'd7;
      34: stateTransition = 11'd7;
      35: stateTransition = 11'd7;
      36: stateTransition = 11'd7;
      37: stateTransition = 11'd7;
      38: stateTransition = 11'd7;
      39: stateTransition = 11'd7;
      40: stateTransition = 11'd7;
      default: stateTransition = 11'bX;
    endcase
    61: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    62: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd21;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd21;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd21;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd21;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd125;
      16: stateTransition = 11'd21;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd21;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd21;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd21;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd21;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd21;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    63: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd55;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    64: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd20;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd20;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd20;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd20;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    65: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd20;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd20;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd20;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd20;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    66: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd76;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd76;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd76;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd51;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd76;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    67: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd44;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd44;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd44;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    68: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd43;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd43;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd43;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd43;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    69: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    70: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd43;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd43;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd43;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd43;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    71: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd46;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd46;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd46;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd46;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    72: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd49;
      17: stateTransition = 11'd48;
      18: stateTransition = 11'd49;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd49;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd49;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    73: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd52;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd52;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd52;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd51;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd52;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    74: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd444;
      2: stateTransition = 11'd444;
      3: stateTransition = 11'd444;
      4: stateTransition = 11'd444;
      5: stateTransition = 11'd444;
      6: stateTransition = 11'd448;
      7: stateTransition = 11'd444;
      8: stateTransition = 11'd444;
      9: stateTransition = 11'd444;
      10: stateTransition = 11'd444;
      11: stateTransition = 11'd444;
      12: stateTransition = 11'd444;
      13: stateTransition = 11'd444;
      14: stateTransition = 11'd444;
      15: stateTransition = 11'd444;
      16: stateTransition = 11'd444;
      17: stateTransition = 11'd444;
      18: stateTransition = 11'd444;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd444;
      22: stateTransition = 11'd444;
      23: stateTransition = 11'd444;
      24: stateTransition = 11'd444;
      25: stateTransition = 11'd444;
      26: stateTransition = 11'd444;
      27: stateTransition = 11'd444;
      28: stateTransition = 11'd444;
      29: stateTransition = 11'd444;
      30: stateTransition = 11'd444;
      31: stateTransition = 11'd444;
      32: stateTransition = 11'd444;
      33: stateTransition = 11'd444;
      34: stateTransition = 11'd444;
      35: stateTransition = 11'd444;
      36: stateTransition = 11'd444;
      37: stateTransition = 11'd444;
      38: stateTransition = 11'd444;
      39: stateTransition = 11'd444;
      40: stateTransition = 11'd444;
      default: stateTransition = 11'bX;
    endcase
    75: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd181;
      2: stateTransition = 11'd181;
      3: stateTransition = 11'd181;
      4: stateTransition = 11'd181;
      5: stateTransition = 11'd181;
      6: stateTransition = 11'd181;
      7: stateTransition = 11'd181;
      8: stateTransition = 11'd133;
      9: stateTransition = 11'd181;
      10: stateTransition = 11'd181;
      11: stateTransition = 11'd181;
      12: stateTransition = 11'd181;
      13: stateTransition = 11'd181;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd181;
      16: stateTransition = 11'd181;
      17: stateTransition = 11'd181;
      18: stateTransition = 11'd181;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd181;
      22: stateTransition = 11'd181;
      23: stateTransition = 11'd181;
      24: stateTransition = 11'd181;
      25: stateTransition = 11'd181;
      26: stateTransition = 11'd181;
      27: stateTransition = 11'd181;
      28: stateTransition = 11'd181;
      29: stateTransition = 11'd181;
      30: stateTransition = 11'd181;
      31: stateTransition = 11'd181;
      32: stateTransition = 11'd181;
      33: stateTransition = 11'd181;
      34: stateTransition = 11'd181;
      35: stateTransition = 11'd181;
      36: stateTransition = 11'd181;
      37: stateTransition = 11'd181;
      38: stateTransition = 11'd181;
      39: stateTransition = 11'd181;
      40: stateTransition = 11'd181;
      default: stateTransition = 11'bX;
    endcase
    76: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd56;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    77: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd16;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd16;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd16;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd16;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    78: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd52;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd52;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd52;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd51;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd52;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    79: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd47;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd47;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd47;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    80: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd74;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd74;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd74;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd74;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    81: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd48;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    82: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd458;
      2: stateTransition = 11'd458;
      3: stateTransition = 11'd458;
      4: stateTransition = 11'd458;
      5: stateTransition = 11'd458;
      6: stateTransition = 11'd458;
      7: stateTransition = 11'd458;
      8: stateTransition = 11'd458;
      9: stateTransition = 11'd458;
      10: stateTransition = 11'd458;
      11: stateTransition = 11'd458;
      12: stateTransition = 11'd458;
      13: stateTransition = 11'd458;
      14: stateTransition = 11'd458;
      15: stateTransition = 11'd9;
      16: stateTransition = 11'd458;
      17: stateTransition = 11'd458;
      18: stateTransition = 11'd458;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd458;
      22: stateTransition = 11'd458;
      23: stateTransition = 11'd458;
      24: stateTransition = 11'd458;
      25: stateTransition = 11'd458;
      26: stateTransition = 11'd458;
      27: stateTransition = 11'd458;
      28: stateTransition = 11'd458;
      29: stateTransition = 11'd458;
      30: stateTransition = 11'd458;
      31: stateTransition = 11'd458;
      32: stateTransition = 11'd458;
      33: stateTransition = 11'd458;
      34: stateTransition = 11'd458;
      35: stateTransition = 11'd458;
      36: stateTransition = 11'd458;
      37: stateTransition = 11'd458;
      38: stateTransition = 11'd458;
      39: stateTransition = 11'd458;
      40: stateTransition = 11'd458;
      default: stateTransition = 11'bX;
    endcase
    83: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd57;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    84: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd50;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd50;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    85: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd46;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd46;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd46;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd46;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    86: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd458;
      2: stateTransition = 11'd458;
      3: stateTransition = 11'd458;
      4: stateTransition = 11'd458;
      5: stateTransition = 11'd458;
      6: stateTransition = 11'd458;
      7: stateTransition = 11'd458;
      8: stateTransition = 11'd458;
      9: stateTransition = 11'd458;
      10: stateTransition = 11'd458;
      11: stateTransition = 11'd458;
      12: stateTransition = 11'd458;
      13: stateTransition = 11'd458;
      14: stateTransition = 11'd458;
      15: stateTransition = 11'd458;
      16: stateTransition = 11'd430;
      17: stateTransition = 11'd458;
      18: stateTransition = 11'd430;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd458;
      22: stateTransition = 11'd458;
      23: stateTransition = 11'd458;
      24: stateTransition = 11'd458;
      25: stateTransition = 11'd430;
      26: stateTransition = 11'd458;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd458;
      29: stateTransition = 11'd430;
      30: stateTransition = 11'd458;
      31: stateTransition = 11'd458;
      32: stateTransition = 11'd458;
      33: stateTransition = 11'd458;
      34: stateTransition = 11'd458;
      35: stateTransition = 11'd458;
      36: stateTransition = 11'd458;
      37: stateTransition = 11'd458;
      38: stateTransition = 11'd458;
      39: stateTransition = 11'd458;
      40: stateTransition = 11'd458;
      default: stateTransition = 11'bX;
    endcase
    87: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd58;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    88: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd75;
      17: stateTransition = 11'd48;
      18: stateTransition = 11'd75;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd75;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd75;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    89: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd439;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd439;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd15;
      12: stateTransition = 11'd439;
      13: stateTransition = 11'd439;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd439;
      16: stateTransition = 11'd439;
      17: stateTransition = 11'd439;
      18: stateTransition = 11'd439;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd439;
      22: stateTransition = 11'd439;
      23: stateTransition = 11'd439;
      24: stateTransition = 11'd439;
      25: stateTransition = 11'd439;
      26: stateTransition = 11'd439;
      27: stateTransition = 11'd439;
      28: stateTransition = 11'd439;
      29: stateTransition = 11'd439;
      30: stateTransition = 11'd439;
      31: stateTransition = 11'd439;
      32: stateTransition = 11'd439;
      33: stateTransition = 11'd439;
      34: stateTransition = 11'd439;
      35: stateTransition = 11'd439;
      36: stateTransition = 11'd439;
      37: stateTransition = 11'd439;
      38: stateTransition = 11'd439;
      39: stateTransition = 11'd439;
      40: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    90: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    91: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd36;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd49;
      17: stateTransition = 11'd48;
      18: stateTransition = 11'd49;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd49;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd49;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      32: stateTransition = 11'd0;
      33: stateTransition = 11'd0;
      34: stateTransition = 11'd0;
      35: stateTransition = 11'd0;
      36: stateTransition = 11'd0;
      37: stateTransition = 11'd0;
      38: stateTransition = 11'd0;
      39: stateTransition = 11'd0;
      40: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    92: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd100;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd100;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd100;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd65;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd100;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    93: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd494;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    94: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd175;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd175;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd175;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd175;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    95: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd60;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    96: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd103;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd103;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd21;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd103;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    97: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd474;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    98: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd135;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd135;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd135;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd23;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd135;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    99: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd106;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd106;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd106;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd25;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd106;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    100: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd122;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd122;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd122;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd26;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd122;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    101: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd28;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd28;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd28;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd29;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd28;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    102: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd30;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd30;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd30;
      12: stateTransition = 11'd31;
      13: stateTransition = 11'd30;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd30;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd30;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd30;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd30;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd30;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd30;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    103: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd32;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd32;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd32;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    104: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd71;
      17: stateTransition = 11'd70;
      18: stateTransition = 11'd71;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd71;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd71;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    105: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd33;
      17: stateTransition = 11'd70;
      18: stateTransition = 11'd33;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd33;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd33;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    106: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd84;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd84;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd84;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    107: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd70;
      18: stateTransition = 11'd27;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd27;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd27;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    108: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd89;
      17: stateTransition = 11'd83;
      18: stateTransition = 11'd89;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd89;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd89;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    109: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd72;
      17: stateTransition = 11'd83;
      18: stateTransition = 11'd72;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd72;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd72;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    110: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd92;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd92;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd92;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    111: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd83;
      18: stateTransition = 11'd27;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd27;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd27;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    112: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd95;
      17: stateTransition = 11'd88;
      18: stateTransition = 11'd95;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd95;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd95;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    113: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd85;
      17: stateTransition = 11'd88;
      18: stateTransition = 11'd85;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd85;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd85;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    114: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd69;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd69;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd69;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    115: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd88;
      18: stateTransition = 11'd27;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd27;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd27;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    116: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd82;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd82;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd82;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd34;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd82;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    117: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd35;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd35;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd35;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd34;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd35;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    118: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd27;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd27;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd27;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd34;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd27;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    119: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd140;
      2: stateTransition = 11'd140;
      3: stateTransition = 11'd140;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd140;
      6: stateTransition = 11'd140;
      7: stateTransition = 11'd140;
      8: stateTransition = 11'd140;
      9: stateTransition = 11'd140;
      10: stateTransition = 11'd140;
      11: stateTransition = 11'd140;
      12: stateTransition = 11'd140;
      13: stateTransition = 11'd140;
      14: stateTransition = 11'd140;
      15: stateTransition = 11'd140;
      16: stateTransition = 11'd140;
      17: stateTransition = 11'd140;
      18: stateTransition = 11'd140;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd140;
      22: stateTransition = 11'd140;
      23: stateTransition = 11'd140;
      24: stateTransition = 11'd140;
      25: stateTransition = 11'd140;
      26: stateTransition = 11'd140;
      27: stateTransition = 11'd140;
      28: stateTransition = 11'd140;
      29: stateTransition = 11'd140;
      30: stateTransition = 11'd140;
      31: stateTransition = 11'd140;
      32: stateTransition = 11'd140;
      33: stateTransition = 11'd140;
      34: stateTransition = 11'd140;
      35: stateTransition = 11'd140;
      36: stateTransition = 11'd140;
      37: stateTransition = 11'd140;
      38: stateTransition = 11'd140;
      39: stateTransition = 11'd140;
      40: stateTransition = 11'd140;
      default: stateTransition = 11'bX;
    endcase
    120: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd105;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd105;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd105;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    121: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    122: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd27;
      2: stateTransition = 11'd27;
      3: stateTransition = 11'd27;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd27;
      8: stateTransition = 11'd27;
      9: stateTransition = 11'd27;
      10: stateTransition = 11'd27;
      11: stateTransition = 11'd27;
      12: stateTransition = 11'd27;
      13: stateTransition = 11'd27;
      14: stateTransition = 11'd27;
      15: stateTransition = 11'd27;
      16: stateTransition = 11'd81;
      17: stateTransition = 11'd27;
      18: stateTransition = 11'd81;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd27;
      22: stateTransition = 11'd27;
      23: stateTransition = 11'd27;
      24: stateTransition = 11'd27;
      25: stateTransition = 11'd81;
      26: stateTransition = 11'd27;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd27;
      29: stateTransition = 11'd81;
      30: stateTransition = 11'd27;
      31: stateTransition = 11'd27;
      32: stateTransition = 11'd27;
      33: stateTransition = 11'd27;
      34: stateTransition = 11'd27;
      35: stateTransition = 11'd27;
      36: stateTransition = 11'd27;
      37: stateTransition = 11'd27;
      38: stateTransition = 11'd27;
      39: stateTransition = 11'd27;
      40: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    123: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd65;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd65;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd65;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd65;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd169;
      16: stateTransition = 11'd65;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd65;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd65;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd65;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd65;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd65;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    124: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd66;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    125: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd149;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    126: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd130;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    127: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd131;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    128: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd465;
      2: stateTransition = 11'd465;
      3: stateTransition = 11'd465;
      4: stateTransition = 11'd465;
      5: stateTransition = 11'd465;
      6: stateTransition = 11'd465;
      7: stateTransition = 11'd465;
      8: stateTransition = 11'd465;
      9: stateTransition = 11'd465;
      10: stateTransition = 11'd465;
      11: stateTransition = 11'd465;
      12: stateTransition = 11'd86;
      13: stateTransition = 11'd465;
      14: stateTransition = 11'd465;
      15: stateTransition = 11'd465;
      16: stateTransition = 11'd465;
      17: stateTransition = 11'd465;
      18: stateTransition = 11'd465;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd465;
      22: stateTransition = 11'd465;
      23: stateTransition = 11'd465;
      24: stateTransition = 11'd465;
      25: stateTransition = 11'd465;
      26: stateTransition = 11'd465;
      27: stateTransition = 11'd465;
      28: stateTransition = 11'd465;
      29: stateTransition = 11'd465;
      30: stateTransition = 11'd465;
      31: stateTransition = 11'd465;
      32: stateTransition = 11'd465;
      33: stateTransition = 11'd465;
      34: stateTransition = 11'd465;
      35: stateTransition = 11'd465;
      36: stateTransition = 11'd465;
      37: stateTransition = 11'd465;
      38: stateTransition = 11'd465;
      39: stateTransition = 11'd465;
      40: stateTransition = 11'd465;
      default: stateTransition = 11'bX;
    endcase
    129: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd96;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd96;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd96;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd128;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd96;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    130: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd123;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd123;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd123;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd26;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd123;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    131: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd140;
      2: stateTransition = 11'd140;
      3: stateTransition = 11'd140;
      4: stateTransition = 11'd140;
      5: stateTransition = 11'd140;
      6: stateTransition = 11'd140;
      7: stateTransition = 11'd178;
      8: stateTransition = 11'd140;
      9: stateTransition = 11'd140;
      10: stateTransition = 11'd140;
      11: stateTransition = 11'd140;
      12: stateTransition = 11'd140;
      13: stateTransition = 11'd140;
      14: stateTransition = 11'd140;
      15: stateTransition = 11'd140;
      16: stateTransition = 11'd140;
      17: stateTransition = 11'd140;
      18: stateTransition = 11'd140;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd140;
      22: stateTransition = 11'd140;
      23: stateTransition = 11'd140;
      24: stateTransition = 11'd140;
      25: stateTransition = 11'd140;
      26: stateTransition = 11'd140;
      27: stateTransition = 11'd140;
      28: stateTransition = 11'd140;
      29: stateTransition = 11'd140;
      30: stateTransition = 11'd140;
      31: stateTransition = 11'd140;
      32: stateTransition = 11'd140;
      33: stateTransition = 11'd140;
      34: stateTransition = 11'd140;
      35: stateTransition = 11'd140;
      36: stateTransition = 11'd140;
      37: stateTransition = 11'd140;
      38: stateTransition = 11'd140;
      39: stateTransition = 11'd140;
      40: stateTransition = 11'd140;
      default: stateTransition = 11'bX;
    endcase
    132: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd80;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd80;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd80;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd80;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    133: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd465;
      2: stateTransition = 11'd465;
      3: stateTransition = 11'd465;
      4: stateTransition = 11'd465;
      5: stateTransition = 11'd465;
      6: stateTransition = 11'd465;
      7: stateTransition = 11'd465;
      8: stateTransition = 11'd465;
      9: stateTransition = 11'd465;
      10: stateTransition = 11'd465;
      11: stateTransition = 11'd465;
      12: stateTransition = 11'd90;
      13: stateTransition = 11'd465;
      14: stateTransition = 11'd465;
      15: stateTransition = 11'd465;
      16: stateTransition = 11'd465;
      17: stateTransition = 11'd465;
      18: stateTransition = 11'd465;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd465;
      22: stateTransition = 11'd465;
      23: stateTransition = 11'd465;
      24: stateTransition = 11'd465;
      25: stateTransition = 11'd465;
      26: stateTransition = 11'd465;
      27: stateTransition = 11'd465;
      28: stateTransition = 11'd465;
      29: stateTransition = 11'd465;
      30: stateTransition = 11'd465;
      31: stateTransition = 11'd465;
      32: stateTransition = 11'd465;
      33: stateTransition = 11'd465;
      34: stateTransition = 11'd465;
      35: stateTransition = 11'd465;
      36: stateTransition = 11'd465;
      37: stateTransition = 11'd465;
      38: stateTransition = 11'd465;
      39: stateTransition = 11'd465;
      40: stateTransition = 11'd465;
      default: stateTransition = 11'bX;
    endcase
    134: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd105;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd105;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd26;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd105;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    135: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd181;
      2: stateTransition = 11'd181;
      3: stateTransition = 11'd181;
      4: stateTransition = 11'd181;
      5: stateTransition = 11'd181;
      6: stateTransition = 11'd181;
      7: stateTransition = 11'd181;
      8: stateTransition = 11'd181;
      9: stateTransition = 11'd181;
      10: stateTransition = 11'd181;
      11: stateTransition = 11'd181;
      12: stateTransition = 11'd181;
      13: stateTransition = 11'd181;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd181;
      16: stateTransition = 11'd181;
      17: stateTransition = 11'd181;
      18: stateTransition = 11'd181;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd181;
      22: stateTransition = 11'd181;
      23: stateTransition = 11'd181;
      24: stateTransition = 11'd181;
      25: stateTransition = 11'd181;
      26: stateTransition = 11'd181;
      27: stateTransition = 11'd181;
      28: stateTransition = 11'd181;
      29: stateTransition = 11'd181;
      30: stateTransition = 11'd181;
      31: stateTransition = 11'd181;
      32: stateTransition = 11'd181;
      33: stateTransition = 11'd181;
      34: stateTransition = 11'd181;
      35: stateTransition = 11'd181;
      36: stateTransition = 11'd181;
      37: stateTransition = 11'd181;
      38: stateTransition = 11'd181;
      39: stateTransition = 11'd181;
      40: stateTransition = 11'd181;
      default: stateTransition = 11'bX;
    endcase
    136: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd132;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    137: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd465;
      2: stateTransition = 11'd465;
      3: stateTransition = 11'd465;
      4: stateTransition = 11'd465;
      5: stateTransition = 11'd465;
      6: stateTransition = 11'd465;
      7: stateTransition = 11'd452;
      8: stateTransition = 11'd465;
      9: stateTransition = 11'd465;
      10: stateTransition = 11'd465;
      11: stateTransition = 11'd465;
      12: stateTransition = 11'd465;
      13: stateTransition = 11'd465;
      14: stateTransition = 11'd465;
      15: stateTransition = 11'd465;
      16: stateTransition = 11'd465;
      17: stateTransition = 11'd465;
      18: stateTransition = 11'd465;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd465;
      22: stateTransition = 11'd465;
      23: stateTransition = 11'd465;
      24: stateTransition = 11'd465;
      25: stateTransition = 11'd465;
      26: stateTransition = 11'd465;
      27: stateTransition = 11'd465;
      28: stateTransition = 11'd465;
      29: stateTransition = 11'd465;
      30: stateTransition = 11'd465;
      31: stateTransition = 11'd465;
      32: stateTransition = 11'd465;
      33: stateTransition = 11'd465;
      34: stateTransition = 11'd465;
      35: stateTransition = 11'd465;
      36: stateTransition = 11'd465;
      37: stateTransition = 11'd465;
      38: stateTransition = 11'd465;
      39: stateTransition = 11'd465;
      40: stateTransition = 11'd465;
      default: stateTransition = 11'bX;
    endcase
    138: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd87;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    139: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd460;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd460;
      10: stateTransition = 11'd93;
      11: stateTransition = 11'd460;
      12: stateTransition = 11'd460;
      13: stateTransition = 11'd460;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd460;
      16: stateTransition = 11'd460;
      17: stateTransition = 11'd460;
      18: stateTransition = 11'd460;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd460;
      22: stateTransition = 11'd460;
      23: stateTransition = 11'd460;
      24: stateTransition = 11'd460;
      25: stateTransition = 11'd460;
      26: stateTransition = 11'd460;
      27: stateTransition = 11'd460;
      28: stateTransition = 11'd460;
      29: stateTransition = 11'd460;
      30: stateTransition = 11'd460;
      31: stateTransition = 11'd460;
      32: stateTransition = 11'd460;
      33: stateTransition = 11'd460;
      34: stateTransition = 11'd460;
      35: stateTransition = 11'd460;
      36: stateTransition = 11'd460;
      37: stateTransition = 11'd460;
      38: stateTransition = 11'd460;
      39: stateTransition = 11'd460;
      40: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    140: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd91;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    141: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd98;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd98;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd98;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    142: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd94;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    143: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd102;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd102;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd102;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    144: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd97;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    145: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd104;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd104;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd104;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    146: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd99;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    147: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd97;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    148: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd107;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd107;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd107;
      12: stateTransition = 11'd108;
      13: stateTransition = 11'd107;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd107;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd107;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd107;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd107;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd107;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd107;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    149: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd101;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    150: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd109;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd109;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd109;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    151: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd110;
      17: stateTransition = 11'd111;
      18: stateTransition = 11'd110;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd110;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd110;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    152: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd111;
      18: stateTransition = 11'd112;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd112;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd112;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    153: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd113;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd113;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd113;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    154: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd111;
      18: stateTransition = 11'd105;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd105;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd105;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    155: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd114;
      17: stateTransition = 11'd115;
      18: stateTransition = 11'd114;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd114;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd114;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    156: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd116;
      17: stateTransition = 11'd115;
      18: stateTransition = 11'd116;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd116;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd116;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    157: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd117;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd117;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd117;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    158: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd115;
      18: stateTransition = 11'd105;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd105;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd105;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    159: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd118;
      17: stateTransition = 11'd119;
      18: stateTransition = 11'd118;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd118;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd118;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    160: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd120;
      17: stateTransition = 11'd119;
      18: stateTransition = 11'd120;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd120;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd120;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    161: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd105;
      18: stateTransition = 11'd121;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd121;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd121;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    162: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd105;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd105;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd105;
      8: stateTransition = 11'd105;
      9: stateTransition = 11'd105;
      10: stateTransition = 11'd105;
      11: stateTransition = 11'd105;
      12: stateTransition = 11'd105;
      13: stateTransition = 11'd105;
      14: stateTransition = 11'd105;
      15: stateTransition = 11'd105;
      16: stateTransition = 11'd105;
      17: stateTransition = 11'd119;
      18: stateTransition = 11'd105;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd105;
      22: stateTransition = 11'd105;
      23: stateTransition = 11'd105;
      24: stateTransition = 11'd105;
      25: stateTransition = 11'd105;
      26: stateTransition = 11'd105;
      27: stateTransition = 11'd105;
      28: stateTransition = 11'd105;
      29: stateTransition = 11'd105;
      30: stateTransition = 11'd105;
      31: stateTransition = 11'd105;
      32: stateTransition = 11'd105;
      33: stateTransition = 11'd105;
      34: stateTransition = 11'd105;
      35: stateTransition = 11'd105;
      36: stateTransition = 11'd105;
      37: stateTransition = 11'd105;
      38: stateTransition = 11'd105;
      39: stateTransition = 11'd105;
      40: stateTransition = 11'd105;
      default: stateTransition = 11'bX;
    endcase
    163: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd152;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd152;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd152;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    164: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    165: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd128;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd128;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd128;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd128;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd206;
      16: stateTransition = 11'd128;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd128;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd128;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd128;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd128;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd128;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    166: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    167: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd181;
      2: stateTransition = 11'd181;
      3: stateTransition = 11'd181;
      4: stateTransition = 11'd181;
      5: stateTransition = 11'd181;
      6: stateTransition = 11'd181;
      7: stateTransition = 11'd181;
      8: stateTransition = 11'd181;
      9: stateTransition = 11'd181;
      10: stateTransition = 11'd181;
      11: stateTransition = 11'd181;
      12: stateTransition = 11'd181;
      13: stateTransition = 11'd181;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd181;
      16: stateTransition = 11'd181;
      17: stateTransition = 11'd181;
      18: stateTransition = 11'd181;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd181;
      22: stateTransition = 11'd181;
      23: stateTransition = 11'd181;
      24: stateTransition = 11'd181;
      25: stateTransition = 11'd181;
      26: stateTransition = 11'd181;
      27: stateTransition = 11'd181;
      28: stateTransition = 11'd181;
      29: stateTransition = 11'd181;
      30: stateTransition = 11'd181;
      31: stateTransition = 11'd181;
      32: stateTransition = 11'd181;
      33: stateTransition = 11'd181;
      34: stateTransition = 11'd181;
      35: stateTransition = 11'd181;
      36: stateTransition = 11'd181;
      37: stateTransition = 11'd181;
      38: stateTransition = 11'd138;
      39: stateTransition = 11'd181;
      40: stateTransition = 11'd181;
      default: stateTransition = 11'bX;
    endcase
    168: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd134;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd134;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd134;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd171;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd134;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    169: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd139;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd139;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd139;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd23;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd139;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    170: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd468;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd468;
      10: stateTransition = 11'd144;
      11: stateTransition = 11'd468;
      12: stateTransition = 11'd468;
      13: stateTransition = 11'd468;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd468;
      16: stateTransition = 11'd468;
      17: stateTransition = 11'd468;
      18: stateTransition = 11'd468;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd468;
      22: stateTransition = 11'd468;
      23: stateTransition = 11'd468;
      24: stateTransition = 11'd468;
      25: stateTransition = 11'd468;
      26: stateTransition = 11'd468;
      27: stateTransition = 11'd468;
      28: stateTransition = 11'd468;
      29: stateTransition = 11'd468;
      30: stateTransition = 11'd468;
      31: stateTransition = 11'd468;
      32: stateTransition = 11'd468;
      33: stateTransition = 11'd468;
      34: stateTransition = 11'd468;
      35: stateTransition = 11'd468;
      36: stateTransition = 11'd468;
      37: stateTransition = 11'd468;
      38: stateTransition = 11'd468;
      39: stateTransition = 11'd468;
      40: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    171: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd137;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    172: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd181;
      2: stateTransition = 11'd181;
      3: stateTransition = 11'd181;
      4: stateTransition = 11'd181;
      5: stateTransition = 11'd181;
      6: stateTransition = 11'd181;
      7: stateTransition = 11'd181;
      8: stateTransition = 11'd181;
      9: stateTransition = 11'd142;
      10: stateTransition = 11'd181;
      11: stateTransition = 11'd181;
      12: stateTransition = 11'd181;
      13: stateTransition = 11'd181;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd181;
      16: stateTransition = 11'd181;
      17: stateTransition = 11'd181;
      18: stateTransition = 11'd181;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd181;
      22: stateTransition = 11'd181;
      23: stateTransition = 11'd181;
      24: stateTransition = 11'd181;
      25: stateTransition = 11'd181;
      26: stateTransition = 11'd181;
      27: stateTransition = 11'd181;
      28: stateTransition = 11'd181;
      29: stateTransition = 11'd181;
      30: stateTransition = 11'd181;
      31: stateTransition = 11'd181;
      32: stateTransition = 11'd181;
      33: stateTransition = 11'd181;
      34: stateTransition = 11'd181;
      35: stateTransition = 11'd181;
      36: stateTransition = 11'd181;
      37: stateTransition = 11'd181;
      38: stateTransition = 11'd181;
      39: stateTransition = 11'd181;
      40: stateTransition = 11'd181;
      default: stateTransition = 11'bX;
    endcase
    173: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd262;
      17: stateTransition = 11'd146;
      18: stateTransition = 11'd262;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd262;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd262;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    174: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd306;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd141;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd185;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd344;
      33: stateTransition = 11'd311;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    175: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd465;
      2: stateTransition = 11'd465;
      3: stateTransition = 11'd465;
      4: stateTransition = 11'd465;
      5: stateTransition = 11'd465;
      6: stateTransition = 11'd465;
      7: stateTransition = 11'd465;
      8: stateTransition = 11'd465;
      9: stateTransition = 11'd465;
      10: stateTransition = 11'd465;
      11: stateTransition = 11'd465;
      12: stateTransition = 11'd465;
      13: stateTransition = 11'd465;
      14: stateTransition = 11'd465;
      15: stateTransition = 11'd465;
      16: stateTransition = 11'd465;
      17: stateTransition = 11'd465;
      18: stateTransition = 11'd465;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd465;
      22: stateTransition = 11'd465;
      23: stateTransition = 11'd465;
      24: stateTransition = 11'd465;
      25: stateTransition = 11'd465;
      26: stateTransition = 11'd465;
      27: stateTransition = 11'd465;
      28: stateTransition = 11'd465;
      29: stateTransition = 11'd465;
      30: stateTransition = 11'd465;
      31: stateTransition = 11'd465;
      32: stateTransition = 11'd465;
      33: stateTransition = 11'd465;
      34: stateTransition = 11'd465;
      35: stateTransition = 11'd465;
      36: stateTransition = 11'd465;
      37: stateTransition = 11'd465;
      38: stateTransition = 11'd465;
      39: stateTransition = 11'd465;
      40: stateTransition = 11'd465;
      default: stateTransition = 11'bX;
    endcase
    176: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd218;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd218;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd218;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd218;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    177: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd143;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    178: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd204;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd204;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd204;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd204;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    179: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd143;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    180: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd145;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd686;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    181: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd154;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd154;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd154;
      12: stateTransition = 11'd156;
      13: stateTransition = 11'd154;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd154;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd154;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd154;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd154;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd154;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd154;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    182: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd147;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    183: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd157;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd157;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd157;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    184: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd158;
      17: stateTransition = 11'd159;
      18: stateTransition = 11'd158;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd158;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd158;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    185: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd151;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    186: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd160;
      17: stateTransition = 11'd159;
      18: stateTransition = 11'd160;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd160;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd160;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    187: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd153;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    188: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd161;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd161;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd161;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    189: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd686;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd155;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    190: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd159;
      18: stateTransition = 11'd152;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd152;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd152;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    191: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd162;
      17: stateTransition = 11'd163;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd162;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd162;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    192: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd164;
      17: stateTransition = 11'd163;
      18: stateTransition = 11'd164;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd164;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd164;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    193: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd152;
      18: stateTransition = 11'd165;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd165;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd165;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    194: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd163;
      18: stateTransition = 11'd152;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd152;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd152;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    195: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd166;
      17: stateTransition = 11'd167;
      18: stateTransition = 11'd166;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd166;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd166;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    196: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd168;
      17: stateTransition = 11'd167;
      18: stateTransition = 11'd168;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd168;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd168;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    197: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd152;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd152;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd152;
      8: stateTransition = 11'd152;
      9: stateTransition = 11'd152;
      10: stateTransition = 11'd152;
      11: stateTransition = 11'd152;
      12: stateTransition = 11'd152;
      13: stateTransition = 11'd152;
      14: stateTransition = 11'd152;
      15: stateTransition = 11'd152;
      16: stateTransition = 11'd152;
      17: stateTransition = 11'd167;
      18: stateTransition = 11'd152;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd152;
      22: stateTransition = 11'd152;
      23: stateTransition = 11'd152;
      24: stateTransition = 11'd152;
      25: stateTransition = 11'd152;
      26: stateTransition = 11'd152;
      27: stateTransition = 11'd152;
      28: stateTransition = 11'd152;
      29: stateTransition = 11'd152;
      30: stateTransition = 11'd152;
      31: stateTransition = 11'd152;
      32: stateTransition = 11'd152;
      33: stateTransition = 11'd152;
      34: stateTransition = 11'd152;
      35: stateTransition = 11'd152;
      36: stateTransition = 11'd152;
      37: stateTransition = 11'd152;
      38: stateTransition = 11'd152;
      39: stateTransition = 11'd152;
      40: stateTransition = 11'd152;
      default: stateTransition = 11'bX;
    endcase
    198: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd186;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd186;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    199: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd170;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    200: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd171;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd171;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd171;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd171;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd251;
      16: stateTransition = 11'd171;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd171;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd171;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd171;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd171;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd171;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    201: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd306;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd277;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd185;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd344;
      33: stateTransition = 11'd311;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    202: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd177;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd177;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd177;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    203: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd210;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    204: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd174;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd174;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd174;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd208;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd174;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    205: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd211;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd592;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    206: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd458;
      2: stateTransition = 11'd458;
      3: stateTransition = 11'd458;
      4: stateTransition = 11'd458;
      5: stateTransition = 11'd458;
      6: stateTransition = 11'd458;
      7: stateTransition = 11'd458;
      8: stateTransition = 11'd458;
      9: stateTransition = 11'd176;
      10: stateTransition = 11'd458;
      11: stateTransition = 11'd458;
      12: stateTransition = 11'd458;
      13: stateTransition = 11'd458;
      14: stateTransition = 11'd458;
      15: stateTransition = 11'd458;
      16: stateTransition = 11'd458;
      17: stateTransition = 11'd458;
      18: stateTransition = 11'd458;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd458;
      22: stateTransition = 11'd458;
      23: stateTransition = 11'd458;
      24: stateTransition = 11'd458;
      25: stateTransition = 11'd458;
      26: stateTransition = 11'd458;
      27: stateTransition = 11'd458;
      28: stateTransition = 11'd458;
      29: stateTransition = 11'd458;
      30: stateTransition = 11'd458;
      31: stateTransition = 11'd458;
      32: stateTransition = 11'd458;
      33: stateTransition = 11'd458;
      34: stateTransition = 11'd458;
      35: stateTransition = 11'd458;
      36: stateTransition = 11'd458;
      37: stateTransition = 11'd458;
      38: stateTransition = 11'd458;
      39: stateTransition = 11'd458;
      40: stateTransition = 11'd458;
      default: stateTransition = 11'bX;
    endcase
    207: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd213;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    208: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd209;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    209: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd465;
      2: stateTransition = 11'd465;
      3: stateTransition = 11'd465;
      4: stateTransition = 11'd465;
      5: stateTransition = 11'd465;
      6: stateTransition = 11'd465;
      7: stateTransition = 11'd465;
      8: stateTransition = 11'd214;
      9: stateTransition = 11'd465;
      10: stateTransition = 11'd465;
      11: stateTransition = 11'd465;
      12: stateTransition = 11'd465;
      13: stateTransition = 11'd465;
      14: stateTransition = 11'd465;
      15: stateTransition = 11'd465;
      16: stateTransition = 11'd465;
      17: stateTransition = 11'd465;
      18: stateTransition = 11'd465;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd465;
      22: stateTransition = 11'd465;
      23: stateTransition = 11'd465;
      24: stateTransition = 11'd465;
      25: stateTransition = 11'd465;
      26: stateTransition = 11'd465;
      27: stateTransition = 11'd465;
      28: stateTransition = 11'd465;
      29: stateTransition = 11'd465;
      30: stateTransition = 11'd465;
      31: stateTransition = 11'd465;
      32: stateTransition = 11'd465;
      33: stateTransition = 11'd465;
      34: stateTransition = 11'd465;
      35: stateTransition = 11'd465;
      36: stateTransition = 11'd465;
      37: stateTransition = 11'd465;
      38: stateTransition = 11'd465;
      39: stateTransition = 11'd465;
      40: stateTransition = 11'd465;
      default: stateTransition = 11'bX;
    endcase
    210: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd205;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd205;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd205;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd205;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    211: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd170;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd215;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    212: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd187;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd480;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    213: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd180;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    214: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd221;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    215: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd222;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    216: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd316;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd179;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd179;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd179;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    217: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd223;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    218: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd150;
      18: stateTransition = 11'd186;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd186;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    219: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd225;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    220: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd189;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    221: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd267;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd271;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd183;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd313;
      33: stateTransition = 11'd275;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    222: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd229;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    223: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd230;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    224: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd182;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd182;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd182;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    225: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd231;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    226: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd233;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    227: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd191;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    228: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd184;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd184;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd184;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    229: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd193;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    230: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd195;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    231: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd188;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd188;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd188;
      12: stateTransition = 11'd190;
      13: stateTransition = 11'd188;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd188;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd188;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd188;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd188;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd188;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd188;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    232: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd197;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    233: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd192;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd192;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd192;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    234: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd194;
      17: stateTransition = 11'd196;
      18: stateTransition = 11'd194;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd194;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd194;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    235: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd198;
      17: stateTransition = 11'd196;
      18: stateTransition = 11'd198;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd198;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd198;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    236: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd199;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd199;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd199;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    237: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd196;
      18: stateTransition = 11'd186;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd186;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    238: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd200;
      17: stateTransition = 11'd201;
      18: stateTransition = 11'd200;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd200;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd200;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    239: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd202;
      17: stateTransition = 11'd201;
      18: stateTransition = 11'd202;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd202;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd202;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    240: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd186;
      18: stateTransition = 11'd203;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd203;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd203;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    241: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd186;
      2: stateTransition = 11'd186;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd186;
      8: stateTransition = 11'd186;
      9: stateTransition = 11'd186;
      10: stateTransition = 11'd186;
      11: stateTransition = 11'd186;
      12: stateTransition = 11'd186;
      13: stateTransition = 11'd186;
      14: stateTransition = 11'd186;
      15: stateTransition = 11'd186;
      16: stateTransition = 11'd186;
      17: stateTransition = 11'd201;
      18: stateTransition = 11'd186;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd186;
      22: stateTransition = 11'd186;
      23: stateTransition = 11'd186;
      24: stateTransition = 11'd186;
      25: stateTransition = 11'd186;
      26: stateTransition = 11'd186;
      27: stateTransition = 11'd186;
      28: stateTransition = 11'd186;
      29: stateTransition = 11'd186;
      30: stateTransition = 11'd186;
      31: stateTransition = 11'd186;
      32: stateTransition = 11'd186;
      33: stateTransition = 11'd186;
      34: stateTransition = 11'd186;
      35: stateTransition = 11'd186;
      36: stateTransition = 11'd186;
      37: stateTransition = 11'd186;
      38: stateTransition = 11'd186;
      39: stateTransition = 11'd186;
      40: stateTransition = 11'd186;
      default: stateTransition = 11'bX;
    endcase
    242: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd238;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd238;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd238;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    243: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd207;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd207;
      9: stateTransition = 11'd207;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd207;
      13: stateTransition = 11'd576;
      14: stateTransition = 11'd207;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd207;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd207;
      22: stateTransition = 11'd207;
      23: stateTransition = 11'd207;
      24: stateTransition = 11'd207;
      25: stateTransition = 11'd207;
      26: stateTransition = 11'd207;
      27: stateTransition = 11'd207;
      28: stateTransition = 11'd207;
      29: stateTransition = 11'd207;
      30: stateTransition = 11'd207;
      31: stateTransition = 11'd207;
      32: stateTransition = 11'd207;
      33: stateTransition = 11'd207;
      34: stateTransition = 11'd207;
      35: stateTransition = 11'd207;
      36: stateTransition = 11'd207;
      37: stateTransition = 11'd207;
      38: stateTransition = 11'd207;
      39: stateTransition = 11'd207;
      40: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    244: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd208;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd208;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd208;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd208;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd291;
      16: stateTransition = 11'd208;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd208;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd208;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd208;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd208;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd208;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    245: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd209;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    246: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd216;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    247: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd255;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    248: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd212;
      17: stateTransition = 11'd358;
      18: stateTransition = 11'd212;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd212;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd253;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd212;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    249: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd256;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    250: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd341;
      17: stateTransition = 11'd224;
      18: stateTransition = 11'd341;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd341;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd341;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    251: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd258;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    252: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd254;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    253: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd226;
      17: stateTransition = 11'd148;
      18: stateTransition = 11'd226;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd226;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd226;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    254: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd260;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    255: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd219;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd545;
      9: stateTransition = 11'd207;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd207;
      13: stateTransition = 11'd576;
      14: stateTransition = 11'd207;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd207;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd207;
      22: stateTransition = 11'd207;
      23: stateTransition = 11'd207;
      24: stateTransition = 11'd207;
      25: stateTransition = 11'd207;
      26: stateTransition = 11'd207;
      27: stateTransition = 11'd207;
      28: stateTransition = 11'd207;
      29: stateTransition = 11'd207;
      30: stateTransition = 11'd207;
      31: stateTransition = 11'd207;
      32: stateTransition = 11'd207;
      33: stateTransition = 11'd207;
      34: stateTransition = 11'd207;
      35: stateTransition = 11'd207;
      36: stateTransition = 11'd207;
      37: stateTransition = 11'd207;
      38: stateTransition = 11'd207;
      39: stateTransition = 11'd207;
      40: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    256: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd220;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd228;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    257: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd304;
      17: stateTransition = 11'd232;
      18: stateTransition = 11'd304;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd304;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd304;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    258: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd265;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd414;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    259: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd263;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    260: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd235;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    261: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd289;
      17: stateTransition = 11'd236;
      18: stateTransition = 11'd289;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd289;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd289;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    262: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd269;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    263: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd227;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    264: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd687;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    265: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd273;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    266: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd234;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    267: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd269;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    268: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd240;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd240;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd240;
      12: stateTransition = 11'd242;
      13: stateTransition = 11'd240;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd240;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd240;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd240;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd240;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd240;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd240;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    269: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd237;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    270: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd243;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd243;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd243;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    271: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd239;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    272: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd244;
      17: stateTransition = 11'd245;
      18: stateTransition = 11'd244;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd244;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd244;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    273: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd484;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    274: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd246;
      17: stateTransition = 11'd245;
      18: stateTransition = 11'd246;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd246;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd246;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    275: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd241;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    276: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd238;
      18: stateTransition = 11'd247;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd247;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd247;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    277: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd245;
      18: stateTransition = 11'd238;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd238;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd238;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    278: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd248;
      17: stateTransition = 11'd249;
      18: stateTransition = 11'd248;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd248;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd248;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    279: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd250;
      17: stateTransition = 11'd249;
      18: stateTransition = 11'd250;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd250;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd250;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    280: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd238;
      2: stateTransition = 11'd238;
      3: stateTransition = 11'd238;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd238;
      8: stateTransition = 11'd238;
      9: stateTransition = 11'd238;
      10: stateTransition = 11'd238;
      11: stateTransition = 11'd238;
      12: stateTransition = 11'd238;
      13: stateTransition = 11'd238;
      14: stateTransition = 11'd238;
      15: stateTransition = 11'd238;
      16: stateTransition = 11'd238;
      17: stateTransition = 11'd249;
      18: stateTransition = 11'd238;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd238;
      22: stateTransition = 11'd238;
      23: stateTransition = 11'd238;
      24: stateTransition = 11'd238;
      25: stateTransition = 11'd238;
      26: stateTransition = 11'd238;
      27: stateTransition = 11'd238;
      28: stateTransition = 11'd238;
      29: stateTransition = 11'd238;
      30: stateTransition = 11'd238;
      31: stateTransition = 11'd238;
      32: stateTransition = 11'd238;
      33: stateTransition = 11'd238;
      34: stateTransition = 11'd238;
      35: stateTransition = 11'd238;
      36: stateTransition = 11'd238;
      37: stateTransition = 11'd238;
      38: stateTransition = 11'd238;
      39: stateTransition = 11'd238;
      40: stateTransition = 11'd238;
      default: stateTransition = 11'bX;
    endcase
    281: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd274;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd274;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd274;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    282: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd252;
      2: stateTransition = 11'd252;
      3: stateTransition = 11'd252;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd252;
      8: stateTransition = 11'd252;
      9: stateTransition = 11'd252;
      10: stateTransition = 11'd252;
      11: stateTransition = 11'd252;
      12: stateTransition = 11'd252;
      13: stateTransition = 11'd567;
      14: stateTransition = 11'd252;
      15: stateTransition = 11'd252;
      16: stateTransition = 11'd252;
      17: stateTransition = 11'd252;
      18: stateTransition = 11'd252;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd252;
      22: stateTransition = 11'd252;
      23: stateTransition = 11'd252;
      24: stateTransition = 11'd252;
      25: stateTransition = 11'd252;
      26: stateTransition = 11'd252;
      27: stateTransition = 11'd252;
      28: stateTransition = 11'd252;
      29: stateTransition = 11'd252;
      30: stateTransition = 11'd252;
      31: stateTransition = 11'd252;
      32: stateTransition = 11'd252;
      33: stateTransition = 11'd252;
      34: stateTransition = 11'd252;
      35: stateTransition = 11'd252;
      36: stateTransition = 11'd252;
      37: stateTransition = 11'd252;
      38: stateTransition = 11'd252;
      39: stateTransition = 11'd252;
      40: stateTransition = 11'd252;
      default: stateTransition = 11'bX;
    endcase
    283: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd253;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd253;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd253;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd253;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd328;
      16: stateTransition = 11'd253;
      17: stateTransition = 11'd358;
      18: stateTransition = 11'd253;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd253;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd253;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd253;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd253;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    284: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd254;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    285: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd261;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    286: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd295;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    287: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd257;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd257;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd257;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd293;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd257;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd393;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    288: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd296;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    289: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd393;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd259;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd259;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd259;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd393;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    290: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd298;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    291: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd294;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    292: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd300;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    293: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd302;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    294: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd290;
      17: stateTransition = 11'd236;
      18: stateTransition = 11'd290;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd290;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd290;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    295: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd252;
      2: stateTransition = 11'd264;
      3: stateTransition = 11'd252;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd252;
      8: stateTransition = 11'd252;
      9: stateTransition = 11'd252;
      10: stateTransition = 11'd252;
      11: stateTransition = 11'd252;
      12: stateTransition = 11'd252;
      13: stateTransition = 11'd567;
      14: stateTransition = 11'd252;
      15: stateTransition = 11'd252;
      16: stateTransition = 11'd252;
      17: stateTransition = 11'd252;
      18: stateTransition = 11'd252;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd252;
      22: stateTransition = 11'd252;
      23: stateTransition = 11'd252;
      24: stateTransition = 11'd252;
      25: stateTransition = 11'd252;
      26: stateTransition = 11'd252;
      27: stateTransition = 11'd252;
      28: stateTransition = 11'd252;
      29: stateTransition = 11'd252;
      30: stateTransition = 11'd252;
      31: stateTransition = 11'd252;
      32: stateTransition = 11'd252;
      33: stateTransition = 11'd252;
      34: stateTransition = 11'd252;
      35: stateTransition = 11'd252;
      36: stateTransition = 11'd252;
      37: stateTransition = 11'd252;
      38: stateTransition = 11'd252;
      39: stateTransition = 11'd252;
      40: stateTransition = 11'd252;
      default: stateTransition = 11'bX;
    endcase
    296: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd265;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd414;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    297: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd358;
      17: stateTransition = 11'd358;
      18: stateTransition = 11'd266;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd266;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd266;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    298: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd315;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd480;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    299: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      17: stateTransition = 11'd236;
      18: stateTransition = 11'd274;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd274;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd274;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    300: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd303;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    301: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd273;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    302: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd316;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd270;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd270;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd270;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    303: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd318;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    304: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd268;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    305: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd279;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    306: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd272;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    307: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd281;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    308: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd278;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd278;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd278;
      12: stateTransition = 11'd280;
      13: stateTransition = 11'd278;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd278;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd278;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd278;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd278;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd278;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd278;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    309: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd276;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    310: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd283;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    311: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd282;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd282;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd282;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    312: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd285;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    313: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd284;
      17: stateTransition = 11'd286;
      18: stateTransition = 11'd284;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd284;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd284;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    314: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd287;
      17: stateTransition = 11'd286;
      18: stateTransition = 11'd287;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd287;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd287;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    315: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      17: stateTransition = 11'd274;
      18: stateTransition = 11'd288;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd288;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd288;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    316: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd274;
      2: stateTransition = 11'd274;
      3: stateTransition = 11'd274;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd274;
      8: stateTransition = 11'd274;
      9: stateTransition = 11'd274;
      10: stateTransition = 11'd274;
      11: stateTransition = 11'd274;
      12: stateTransition = 11'd274;
      13: stateTransition = 11'd274;
      14: stateTransition = 11'd274;
      15: stateTransition = 11'd274;
      16: stateTransition = 11'd274;
      17: stateTransition = 11'd286;
      18: stateTransition = 11'd274;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd274;
      22: stateTransition = 11'd274;
      23: stateTransition = 11'd274;
      24: stateTransition = 11'd274;
      25: stateTransition = 11'd274;
      26: stateTransition = 11'd274;
      27: stateTransition = 11'd274;
      28: stateTransition = 11'd274;
      29: stateTransition = 11'd274;
      30: stateTransition = 11'd274;
      31: stateTransition = 11'd274;
      32: stateTransition = 11'd274;
      33: stateTransition = 11'd274;
      34: stateTransition = 11'd274;
      35: stateTransition = 11'd274;
      36: stateTransition = 11'd274;
      37: stateTransition = 11'd274;
      38: stateTransition = 11'd274;
      39: stateTransition = 11'd274;
      40: stateTransition = 11'd274;
      default: stateTransition = 11'bX;
    endcase
    317: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd316;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd316;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd316;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd316;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    318: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd292;
      2: stateTransition = 11'd292;
      3: stateTransition = 11'd292;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd292;
      8: stateTransition = 11'd292;
      9: stateTransition = 11'd292;
      10: stateTransition = 11'd292;
      11: stateTransition = 11'd292;
      12: stateTransition = 11'd292;
      13: stateTransition = 11'd558;
      14: stateTransition = 11'd292;
      15: stateTransition = 11'd292;
      16: stateTransition = 11'd292;
      17: stateTransition = 11'd292;
      18: stateTransition = 11'd292;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd292;
      22: stateTransition = 11'd292;
      23: stateTransition = 11'd292;
      24: stateTransition = 11'd292;
      25: stateTransition = 11'd292;
      26: stateTransition = 11'd292;
      27: stateTransition = 11'd292;
      28: stateTransition = 11'd292;
      29: stateTransition = 11'd292;
      30: stateTransition = 11'd292;
      31: stateTransition = 11'd292;
      32: stateTransition = 11'd292;
      33: stateTransition = 11'd292;
      34: stateTransition = 11'd292;
      35: stateTransition = 11'd292;
      36: stateTransition = 11'd292;
      37: stateTransition = 11'd292;
      38: stateTransition = 11'd292;
      39: stateTransition = 11'd292;
      40: stateTransition = 11'd292;
      default: stateTransition = 11'bX;
    endcase
    319: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd293;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd293;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd293;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd293;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd368;
      16: stateTransition = 11'd293;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd293;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd293;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd293;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd293;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd293;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    320: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd294;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    321: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd301;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    322: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd332;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    323: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd421;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd421;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd421;
      12: stateTransition = 11'd421;
      13: stateTransition = 11'd421;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd421;
      16: stateTransition = 11'd297;
      17: stateTransition = 11'd421;
      18: stateTransition = 11'd297;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd421;
      22: stateTransition = 11'd421;
      23: stateTransition = 11'd421;
      24: stateTransition = 11'd421;
      25: stateTransition = 11'd297;
      26: stateTransition = 11'd421;
      27: stateTransition = 11'd330;
      28: stateTransition = 11'd421;
      29: stateTransition = 11'd297;
      30: stateTransition = 11'd421;
      31: stateTransition = 11'd421;
      32: stateTransition = 11'd421;
      33: stateTransition = 11'd421;
      34: stateTransition = 11'd421;
      35: stateTransition = 11'd421;
      36: stateTransition = 11'd421;
      37: stateTransition = 11'd421;
      38: stateTransition = 11'd421;
      39: stateTransition = 11'd421;
      40: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    324: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd333;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    325: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd421;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd421;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd421;
      12: stateTransition = 11'd421;
      13: stateTransition = 11'd421;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd421;
      16: stateTransition = 11'd412;
      17: stateTransition = 11'd299;
      18: stateTransition = 11'd412;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd421;
      22: stateTransition = 11'd421;
      23: stateTransition = 11'd421;
      24: stateTransition = 11'd421;
      25: stateTransition = 11'd412;
      26: stateTransition = 11'd421;
      27: stateTransition = 11'd421;
      28: stateTransition = 11'd421;
      29: stateTransition = 11'd412;
      30: stateTransition = 11'd421;
      31: stateTransition = 11'd421;
      32: stateTransition = 11'd421;
      33: stateTransition = 11'd421;
      34: stateTransition = 11'd421;
      35: stateTransition = 11'd421;
      36: stateTransition = 11'd421;
      37: stateTransition = 11'd421;
      38: stateTransition = 11'd421;
      39: stateTransition = 11'd421;
      40: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    326: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd335;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    327: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd331;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    328: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd337;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    329: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd339;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    330: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd309;
      17: stateTransition = 11'd232;
      18: stateTransition = 11'd309;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd309;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd309;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    331: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd340;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    332: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd292;
      2: stateTransition = 11'd292;
      3: stateTransition = 11'd292;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd292;
      8: stateTransition = 11'd292;
      9: stateTransition = 11'd292;
      10: stateTransition = 11'd292;
      11: stateTransition = 11'd292;
      12: stateTransition = 11'd292;
      13: stateTransition = 11'd558;
      14: stateTransition = 11'd305;
      15: stateTransition = 11'd292;
      16: stateTransition = 11'd292;
      17: stateTransition = 11'd292;
      18: stateTransition = 11'd292;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd292;
      22: stateTransition = 11'd292;
      23: stateTransition = 11'd292;
      24: stateTransition = 11'd292;
      25: stateTransition = 11'd292;
      26: stateTransition = 11'd292;
      27: stateTransition = 11'd292;
      28: stateTransition = 11'd292;
      29: stateTransition = 11'd292;
      30: stateTransition = 11'd292;
      31: stateTransition = 11'd292;
      32: stateTransition = 11'd292;
      33: stateTransition = 11'd292;
      34: stateTransition = 11'd292;
      35: stateTransition = 11'd292;
      36: stateTransition = 11'd292;
      37: stateTransition = 11'd292;
      38: stateTransition = 11'd292;
      39: stateTransition = 11'd292;
      40: stateTransition = 11'd292;
      default: stateTransition = 11'bX;
    endcase
    333: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd318;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    334: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd308;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    335: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd345;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    336: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd346;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    337: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd384;
      17: stateTransition = 11'd307;
      18: stateTransition = 11'd384;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd384;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd384;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd393;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    338: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd347;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    339: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd349;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    340: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd350;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    341: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd351;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    342: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd342;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    343: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd321;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    344: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd366;
      17: stateTransition = 11'd312;
      18: stateTransition = 11'd366;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd366;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd366;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    345: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd310;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    346: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd323;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    347: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd314;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    348: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd319;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd319;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd319;
      12: stateTransition = 11'd322;
      13: stateTransition = 11'd319;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd319;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd319;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd319;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd319;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd319;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd319;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    349: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd317;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    350: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd316;
      17: stateTransition = 11'd316;
      18: stateTransition = 11'd324;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd324;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd324;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    351: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd352;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    352: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd325;
      17: stateTransition = 11'd326;
      18: stateTransition = 11'd325;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd325;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd325;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    353: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd320;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    354: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd327;
      17: stateTransition = 11'd326;
      18: stateTransition = 11'd327;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd327;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd327;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    355: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd316;
      2: stateTransition = 11'd316;
      3: stateTransition = 11'd316;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd316;
      8: stateTransition = 11'd316;
      9: stateTransition = 11'd316;
      10: stateTransition = 11'd316;
      11: stateTransition = 11'd316;
      12: stateTransition = 11'd316;
      13: stateTransition = 11'd316;
      14: stateTransition = 11'd316;
      15: stateTransition = 11'd316;
      16: stateTransition = 11'd316;
      17: stateTransition = 11'd326;
      18: stateTransition = 11'd316;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd316;
      22: stateTransition = 11'd316;
      23: stateTransition = 11'd316;
      24: stateTransition = 11'd316;
      25: stateTransition = 11'd316;
      26: stateTransition = 11'd316;
      27: stateTransition = 11'd316;
      28: stateTransition = 11'd316;
      29: stateTransition = 11'd316;
      30: stateTransition = 11'd316;
      31: stateTransition = 11'd316;
      32: stateTransition = 11'd316;
      33: stateTransition = 11'd316;
      34: stateTransition = 11'd316;
      35: stateTransition = 11'd316;
      36: stateTransition = 11'd316;
      37: stateTransition = 11'd316;
      38: stateTransition = 11'd316;
      39: stateTransition = 11'd316;
      40: stateTransition = 11'd316;
      default: stateTransition = 11'bX;
    endcase
    356: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd358;
      17: stateTransition = 11'd358;
      18: stateTransition = 11'd358;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd358;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd358;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    357: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    358: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd330;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd330;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd330;
      12: stateTransition = 11'd421;
      13: stateTransition = 11'd330;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd398;
      16: stateTransition = 11'd330;
      17: stateTransition = 11'd421;
      18: stateTransition = 11'd330;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd421;
      22: stateTransition = 11'd421;
      23: stateTransition = 11'd421;
      24: stateTransition = 11'd421;
      25: stateTransition = 11'd330;
      26: stateTransition = 11'd421;
      27: stateTransition = 11'd421;
      28: stateTransition = 11'd421;
      29: stateTransition = 11'd330;
      30: stateTransition = 11'd421;
      31: stateTransition = 11'd421;
      32: stateTransition = 11'd330;
      33: stateTransition = 11'd421;
      34: stateTransition = 11'd421;
      35: stateTransition = 11'd421;
      36: stateTransition = 11'd421;
      37: stateTransition = 11'd421;
      38: stateTransition = 11'd421;
      39: stateTransition = 11'd330;
      40: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    359: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd331;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    360: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd329;
      2: stateTransition = 11'd329;
      3: stateTransition = 11'd329;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd329;
      8: stateTransition = 11'd329;
      9: stateTransition = 11'd329;
      10: stateTransition = 11'd329;
      11: stateTransition = 11'd329;
      12: stateTransition = 11'd329;
      13: stateTransition = 11'd343;
      14: stateTransition = 11'd329;
      15: stateTransition = 11'd329;
      16: stateTransition = 11'd329;
      17: stateTransition = 11'd329;
      18: stateTransition = 11'd329;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd329;
      22: stateTransition = 11'd329;
      23: stateTransition = 11'd329;
      24: stateTransition = 11'd329;
      25: stateTransition = 11'd329;
      26: stateTransition = 11'd329;
      27: stateTransition = 11'd329;
      28: stateTransition = 11'd329;
      29: stateTransition = 11'd329;
      30: stateTransition = 11'd329;
      31: stateTransition = 11'd329;
      32: stateTransition = 11'd329;
      33: stateTransition = 11'd329;
      34: stateTransition = 11'd329;
      35: stateTransition = 11'd329;
      36: stateTransition = 11'd329;
      37: stateTransition = 11'd329;
      38: stateTransition = 11'd329;
      39: stateTransition = 11'd329;
      40: stateTransition = 11'd329;
      default: stateTransition = 11'bX;
    endcase
    361: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd338;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    362: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd373;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    363: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd439;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd439;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd439;
      12: stateTransition = 11'd439;
      13: stateTransition = 11'd439;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd439;
      16: stateTransition = 11'd334;
      17: stateTransition = 11'd439;
      18: stateTransition = 11'd334;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd439;
      22: stateTransition = 11'd439;
      23: stateTransition = 11'd439;
      24: stateTransition = 11'd439;
      25: stateTransition = 11'd334;
      26: stateTransition = 11'd439;
      27: stateTransition = 11'd370;
      28: stateTransition = 11'd439;
      29: stateTransition = 11'd334;
      30: stateTransition = 11'd439;
      31: stateTransition = 11'd439;
      32: stateTransition = 11'd439;
      33: stateTransition = 11'd439;
      34: stateTransition = 11'd439;
      35: stateTransition = 11'd439;
      36: stateTransition = 11'd439;
      37: stateTransition = 11'd439;
      38: stateTransition = 11'd439;
      39: stateTransition = 11'd439;
      40: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    364: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd374;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    365: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd439;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd439;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd439;
      12: stateTransition = 11'd439;
      13: stateTransition = 11'd439;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd439;
      16: stateTransition = 11'd439;
      17: stateTransition = 11'd439;
      18: stateTransition = 11'd336;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd439;
      22: stateTransition = 11'd439;
      23: stateTransition = 11'd439;
      24: stateTransition = 11'd439;
      25: stateTransition = 11'd336;
      26: stateTransition = 11'd439;
      27: stateTransition = 11'd439;
      28: stateTransition = 11'd439;
      29: stateTransition = 11'd336;
      30: stateTransition = 11'd439;
      31: stateTransition = 11'd439;
      32: stateTransition = 11'd439;
      33: stateTransition = 11'd439;
      34: stateTransition = 11'd439;
      35: stateTransition = 11'd439;
      36: stateTransition = 11'd439;
      37: stateTransition = 11'd439;
      38: stateTransition = 11'd439;
      39: stateTransition = 11'd439;
      40: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    366: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd376;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    367: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd371;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    368: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd378;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    369: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd380;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    370: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd381;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    371: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    372: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd367;
      17: stateTransition = 11'd312;
      18: stateTransition = 11'd367;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd367;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd367;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    373: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd356;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    374: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd354;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    375: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd421;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd421;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd421;
      12: stateTransition = 11'd421;
      13: stateTransition = 11'd421;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd421;
      16: stateTransition = 11'd421;
      17: stateTransition = 11'd421;
      18: stateTransition = 11'd348;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd421;
      22: stateTransition = 11'd421;
      23: stateTransition = 11'd421;
      24: stateTransition = 11'd421;
      25: stateTransition = 11'd348;
      26: stateTransition = 11'd421;
      27: stateTransition = 11'd421;
      28: stateTransition = 11'd421;
      29: stateTransition = 11'd348;
      30: stateTransition = 11'd421;
      31: stateTransition = 11'd421;
      32: stateTransition = 11'd421;
      33: stateTransition = 11'd421;
      34: stateTransition = 11'd421;
      35: stateTransition = 11'd421;
      36: stateTransition = 11'd421;
      37: stateTransition = 11'd421;
      38: stateTransition = 11'd421;
      39: stateTransition = 11'd421;
      40: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    376: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd358;
      17: stateTransition = 11'd312;
      18: stateTransition = 11'd358;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd358;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd358;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    377: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd359;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    378: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd357;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    379: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd393;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd355;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd355;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd355;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd393;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    380: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd361;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    381: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd363;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    382: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd360;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd360;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd360;
      12: stateTransition = 11'd362;
      13: stateTransition = 11'd360;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd360;
      17: stateTransition = 11'd358;
      18: stateTransition = 11'd360;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd360;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd360;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd360;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd360;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    383: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd365;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    384: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd358;
      2: stateTransition = 11'd358;
      3: stateTransition = 11'd358;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd358;
      8: stateTransition = 11'd358;
      9: stateTransition = 11'd358;
      10: stateTransition = 11'd358;
      11: stateTransition = 11'd358;
      12: stateTransition = 11'd358;
      13: stateTransition = 11'd358;
      14: stateTransition = 11'd358;
      15: stateTransition = 11'd358;
      16: stateTransition = 11'd358;
      17: stateTransition = 11'd358;
      18: stateTransition = 11'd364;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd358;
      22: stateTransition = 11'd358;
      23: stateTransition = 11'd358;
      24: stateTransition = 11'd358;
      25: stateTransition = 11'd364;
      26: stateTransition = 11'd358;
      27: stateTransition = 11'd358;
      28: stateTransition = 11'd358;
      29: stateTransition = 11'd364;
      30: stateTransition = 11'd358;
      31: stateTransition = 11'd358;
      32: stateTransition = 11'd358;
      33: stateTransition = 11'd358;
      34: stateTransition = 11'd358;
      35: stateTransition = 11'd358;
      36: stateTransition = 11'd358;
      37: stateTransition = 11'd358;
      38: stateTransition = 11'd358;
      39: stateTransition = 11'd358;
      40: stateTransition = 11'd358;
      default: stateTransition = 11'bX;
    endcase
    385: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd393;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd393;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd393;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd393;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd393;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    386: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    387: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd370;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd370;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd370;
      12: stateTransition = 11'd439;
      13: stateTransition = 11'd370;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd424;
      16: stateTransition = 11'd370;
      17: stateTransition = 11'd439;
      18: stateTransition = 11'd370;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd439;
      22: stateTransition = 11'd439;
      23: stateTransition = 11'd439;
      24: stateTransition = 11'd439;
      25: stateTransition = 11'd370;
      26: stateTransition = 11'd439;
      27: stateTransition = 11'd439;
      28: stateTransition = 11'd439;
      29: stateTransition = 11'd370;
      30: stateTransition = 11'd439;
      31: stateTransition = 11'd439;
      32: stateTransition = 11'd370;
      33: stateTransition = 11'd439;
      34: stateTransition = 11'd439;
      35: stateTransition = 11'd439;
      36: stateTransition = 11'd439;
      37: stateTransition = 11'd439;
      38: stateTransition = 11'd439;
      39: stateTransition = 11'd370;
      40: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    388: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd371;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    389: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd379;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    390: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd402;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    391: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd460;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd460;
      10: stateTransition = 11'd460;
      11: stateTransition = 11'd460;
      12: stateTransition = 11'd460;
      13: stateTransition = 11'd460;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd460;
      16: stateTransition = 11'd375;
      17: stateTransition = 11'd460;
      18: stateTransition = 11'd375;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd460;
      22: stateTransition = 11'd460;
      23: stateTransition = 11'd460;
      24: stateTransition = 11'd460;
      25: stateTransition = 11'd375;
      26: stateTransition = 11'd460;
      27: stateTransition = 11'd400;
      28: stateTransition = 11'd460;
      29: stateTransition = 11'd375;
      30: stateTransition = 11'd460;
      31: stateTransition = 11'd460;
      32: stateTransition = 11'd460;
      33: stateTransition = 11'd460;
      34: stateTransition = 11'd460;
      35: stateTransition = 11'd460;
      36: stateTransition = 11'd460;
      37: stateTransition = 11'd460;
      38: stateTransition = 11'd460;
      39: stateTransition = 11'd460;
      40: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    392: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd403;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    393: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd415;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd415;
      10: stateTransition = 11'd460;
      11: stateTransition = 11'd415;
      12: stateTransition = 11'd377;
      13: stateTransition = 11'd415;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd460;
      16: stateTransition = 11'd415;
      17: stateTransition = 11'd460;
      18: stateTransition = 11'd415;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd460;
      22: stateTransition = 11'd460;
      23: stateTransition = 11'd460;
      24: stateTransition = 11'd460;
      25: stateTransition = 11'd415;
      26: stateTransition = 11'd460;
      27: stateTransition = 11'd460;
      28: stateTransition = 11'd460;
      29: stateTransition = 11'd415;
      30: stateTransition = 11'd460;
      31: stateTransition = 11'd460;
      32: stateTransition = 11'd415;
      33: stateTransition = 11'd460;
      34: stateTransition = 11'd460;
      35: stateTransition = 11'd460;
      36: stateTransition = 11'd460;
      37: stateTransition = 11'd460;
      38: stateTransition = 11'd460;
      39: stateTransition = 11'd415;
      40: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    394: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd405;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    395: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    396: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd407;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    397: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd409;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    398: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    399: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd393;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd393;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd393;
      12: stateTransition = 11'd393;
      13: stateTransition = 11'd393;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd388;
      17: stateTransition = 11'd307;
      18: stateTransition = 11'd388;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd388;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd388;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd393;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd393;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    400: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd389;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    401: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd386;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    402: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd418;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd418;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd418;
      12: stateTransition = 11'd387;
      13: stateTransition = 11'd418;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd439;
      16: stateTransition = 11'd418;
      17: stateTransition = 11'd439;
      18: stateTransition = 11'd418;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd439;
      22: stateTransition = 11'd439;
      23: stateTransition = 11'd439;
      24: stateTransition = 11'd439;
      25: stateTransition = 11'd418;
      26: stateTransition = 11'd439;
      27: stateTransition = 11'd439;
      28: stateTransition = 11'd439;
      29: stateTransition = 11'd418;
      30: stateTransition = 11'd439;
      31: stateTransition = 11'd439;
      32: stateTransition = 11'd418;
      33: stateTransition = 11'd439;
      34: stateTransition = 11'd439;
      35: stateTransition = 11'd439;
      36: stateTransition = 11'd439;
      37: stateTransition = 11'd439;
      38: stateTransition = 11'd439;
      39: stateTransition = 11'd418;
      40: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    403: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd392;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    404: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd488;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    405: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd423;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd423;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd423;
      12: stateTransition = 11'd391;
      13: stateTransition = 11'd423;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd421;
      16: stateTransition = 11'd423;
      17: stateTransition = 11'd421;
      18: stateTransition = 11'd423;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd421;
      22: stateTransition = 11'd421;
      23: stateTransition = 11'd421;
      24: stateTransition = 11'd421;
      25: stateTransition = 11'd423;
      26: stateTransition = 11'd421;
      27: stateTransition = 11'd421;
      28: stateTransition = 11'd421;
      29: stateTransition = 11'd423;
      30: stateTransition = 11'd421;
      31: stateTransition = 11'd421;
      32: stateTransition = 11'd423;
      33: stateTransition = 11'd421;
      34: stateTransition = 11'd421;
      35: stateTransition = 11'd421;
      36: stateTransition = 11'd421;
      37: stateTransition = 11'd421;
      38: stateTransition = 11'd421;
      39: stateTransition = 11'd423;
      40: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    406: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd394;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    407: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd390;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    408: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd396;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    409: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd393;
      2: stateTransition = 11'd393;
      3: stateTransition = 11'd395;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd393;
      8: stateTransition = 11'd393;
      9: stateTransition = 11'd395;
      10: stateTransition = 11'd393;
      11: stateTransition = 11'd395;
      12: stateTransition = 11'd397;
      13: stateTransition = 11'd395;
      14: stateTransition = 11'd393;
      15: stateTransition = 11'd393;
      16: stateTransition = 11'd395;
      17: stateTransition = 11'd393;
      18: stateTransition = 11'd395;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd393;
      22: stateTransition = 11'd393;
      23: stateTransition = 11'd393;
      24: stateTransition = 11'd393;
      25: stateTransition = 11'd395;
      26: stateTransition = 11'd393;
      27: stateTransition = 11'd393;
      28: stateTransition = 11'd393;
      29: stateTransition = 11'd395;
      30: stateTransition = 11'd393;
      31: stateTransition = 11'd393;
      32: stateTransition = 11'd395;
      33: stateTransition = 11'd393;
      34: stateTransition = 11'd393;
      35: stateTransition = 11'd393;
      36: stateTransition = 11'd393;
      37: stateTransition = 11'd393;
      38: stateTransition = 11'd393;
      39: stateTransition = 11'd395;
      40: stateTransition = 11'd393;
      default: stateTransition = 11'bX;
    endcase
    410: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd421;
      2: stateTransition = 11'd421;
      3: stateTransition = 11'd421;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd421;
      8: stateTransition = 11'd421;
      9: stateTransition = 11'd421;
      10: stateTransition = 11'd421;
      11: stateTransition = 11'd421;
      12: stateTransition = 11'd421;
      13: stateTransition = 11'd421;
      14: stateTransition = 11'd421;
      15: stateTransition = 11'd421;
      16: stateTransition = 11'd421;
      17: stateTransition = 11'd421;
      18: stateTransition = 11'd421;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd421;
      22: stateTransition = 11'd421;
      23: stateTransition = 11'd421;
      24: stateTransition = 11'd421;
      25: stateTransition = 11'd421;
      26: stateTransition = 11'd421;
      27: stateTransition = 11'd421;
      28: stateTransition = 11'd421;
      29: stateTransition = 11'd421;
      30: stateTransition = 11'd421;
      31: stateTransition = 11'd421;
      32: stateTransition = 11'd421;
      33: stateTransition = 11'd421;
      34: stateTransition = 11'd421;
      35: stateTransition = 11'd421;
      36: stateTransition = 11'd421;
      37: stateTransition = 11'd421;
      38: stateTransition = 11'd421;
      39: stateTransition = 11'd421;
      40: stateTransition = 11'd421;
      default: stateTransition = 11'bX;
    endcase
    411: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd399;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd677;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd399;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd399;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd399;
      35: stateTransition = 11'd399;
      36: stateTransition = 11'd399;
      37: stateTransition = 11'd399;
      38: stateTransition = 11'd399;
      39: stateTransition = 11'd399;
      40: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    412: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd400;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd400;
      10: stateTransition = 11'd460;
      11: stateTransition = 11'd400;
      12: stateTransition = 11'd460;
      13: stateTransition = 11'd400;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd443;
      16: stateTransition = 11'd400;
      17: stateTransition = 11'd460;
      18: stateTransition = 11'd400;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd460;
      22: stateTransition = 11'd460;
      23: stateTransition = 11'd460;
      24: stateTransition = 11'd460;
      25: stateTransition = 11'd400;
      26: stateTransition = 11'd460;
      27: stateTransition = 11'd460;
      28: stateTransition = 11'd460;
      29: stateTransition = 11'd400;
      30: stateTransition = 11'd460;
      31: stateTransition = 11'd460;
      32: stateTransition = 11'd400;
      33: stateTransition = 11'd460;
      34: stateTransition = 11'd460;
      35: stateTransition = 11'd460;
      36: stateTransition = 11'd460;
      37: stateTransition = 11'd460;
      38: stateTransition = 11'd460;
      39: stateTransition = 11'd400;
      40: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    413: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd401;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    414: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd408;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    415: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd428;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    416: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd468;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd468;
      10: stateTransition = 11'd468;
      11: stateTransition = 11'd468;
      12: stateTransition = 11'd468;
      13: stateTransition = 11'd468;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd468;
      16: stateTransition = 11'd404;
      17: stateTransition = 11'd468;
      18: stateTransition = 11'd404;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd468;
      22: stateTransition = 11'd468;
      23: stateTransition = 11'd468;
      24: stateTransition = 11'd468;
      25: stateTransition = 11'd404;
      26: stateTransition = 11'd468;
      27: stateTransition = 11'd426;
      28: stateTransition = 11'd468;
      29: stateTransition = 11'd404;
      30: stateTransition = 11'd468;
      31: stateTransition = 11'd468;
      32: stateTransition = 11'd468;
      33: stateTransition = 11'd468;
      34: stateTransition = 11'd468;
      35: stateTransition = 11'd468;
      36: stateTransition = 11'd468;
      37: stateTransition = 11'd468;
      38: stateTransition = 11'd468;
      39: stateTransition = 11'd468;
      40: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    417: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd429;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    418: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd468;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd468;
      10: stateTransition = 11'd468;
      11: stateTransition = 11'd468;
      12: stateTransition = 11'd406;
      13: stateTransition = 11'd468;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd468;
      16: stateTransition = 11'd468;
      17: stateTransition = 11'd468;
      18: stateTransition = 11'd468;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd468;
      22: stateTransition = 11'd468;
      23: stateTransition = 11'd468;
      24: stateTransition = 11'd468;
      25: stateTransition = 11'd468;
      26: stateTransition = 11'd468;
      27: stateTransition = 11'd468;
      28: stateTransition = 11'd468;
      29: stateTransition = 11'd468;
      30: stateTransition = 11'd468;
      31: stateTransition = 11'd468;
      32: stateTransition = 11'd468;
      33: stateTransition = 11'd468;
      34: stateTransition = 11'd468;
      35: stateTransition = 11'd468;
      36: stateTransition = 11'd468;
      37: stateTransition = 11'd468;
      38: stateTransition = 11'd468;
      39: stateTransition = 11'd468;
      40: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    419: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd431;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    420: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd427;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    421: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd433;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    422: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    423: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd399;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd677;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd399;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd416;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd399;
      35: stateTransition = 11'd399;
      36: stateTransition = 11'd399;
      37: stateTransition = 11'd399;
      38: stateTransition = 11'd399;
      39: stateTransition = 11'd399;
      40: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    424: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd417;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    425: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd399;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd677;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd419;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd399;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd399;
      35: stateTransition = 11'd399;
      36: stateTransition = 11'd399;
      37: stateTransition = 11'd399;
      38: stateTransition = 11'd399;
      39: stateTransition = 11'd399;
      40: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    426: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd420;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    427: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd399;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd422;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd677;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd399;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd399;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd399;
      35: stateTransition = 11'd399;
      36: stateTransition = 11'd399;
      37: stateTransition = 11'd399;
      38: stateTransition = 11'd399;
      39: stateTransition = 11'd399;
      40: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    428: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd439;
      2: stateTransition = 11'd439;
      3: stateTransition = 11'd439;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd439;
      8: stateTransition = 11'd439;
      9: stateTransition = 11'd439;
      10: stateTransition = 11'd439;
      11: stateTransition = 11'd439;
      12: stateTransition = 11'd439;
      13: stateTransition = 11'd439;
      14: stateTransition = 11'd439;
      15: stateTransition = 11'd439;
      16: stateTransition = 11'd439;
      17: stateTransition = 11'd439;
      18: stateTransition = 11'd439;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd439;
      22: stateTransition = 11'd439;
      23: stateTransition = 11'd439;
      24: stateTransition = 11'd439;
      25: stateTransition = 11'd439;
      26: stateTransition = 11'd439;
      27: stateTransition = 11'd439;
      28: stateTransition = 11'd439;
      29: stateTransition = 11'd439;
      30: stateTransition = 11'd439;
      31: stateTransition = 11'd439;
      32: stateTransition = 11'd439;
      33: stateTransition = 11'd439;
      34: stateTransition = 11'd439;
      35: stateTransition = 11'd439;
      36: stateTransition = 11'd439;
      37: stateTransition = 11'd439;
      38: stateTransition = 11'd439;
      39: stateTransition = 11'd439;
      40: stateTransition = 11'd439;
      default: stateTransition = 11'bX;
    endcase
    429: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd460;
      2: stateTransition = 11'd460;
      3: stateTransition = 11'd460;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd443;
      7: stateTransition = 11'd460;
      8: stateTransition = 11'd460;
      9: stateTransition = 11'd460;
      10: stateTransition = 11'd460;
      11: stateTransition = 11'd460;
      12: stateTransition = 11'd460;
      13: stateTransition = 11'd460;
      14: stateTransition = 11'd460;
      15: stateTransition = 11'd460;
      16: stateTransition = 11'd460;
      17: stateTransition = 11'd460;
      18: stateTransition = 11'd460;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd460;
      22: stateTransition = 11'd460;
      23: stateTransition = 11'd460;
      24: stateTransition = 11'd460;
      25: stateTransition = 11'd460;
      26: stateTransition = 11'd460;
      27: stateTransition = 11'd460;
      28: stateTransition = 11'd460;
      29: stateTransition = 11'd460;
      30: stateTransition = 11'd460;
      31: stateTransition = 11'd460;
      32: stateTransition = 11'd460;
      33: stateTransition = 11'd460;
      34: stateTransition = 11'd460;
      35: stateTransition = 11'd460;
      36: stateTransition = 11'd460;
      37: stateTransition = 11'd460;
      38: stateTransition = 11'd460;
      39: stateTransition = 11'd460;
      40: stateTransition = 11'd460;
      default: stateTransition = 11'bX;
    endcase
    430: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd425;
      2: stateTransition = 11'd425;
      3: stateTransition = 11'd425;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd437;
      8: stateTransition = 11'd425;
      9: stateTransition = 11'd425;
      10: stateTransition = 11'd425;
      11: stateTransition = 11'd425;
      12: stateTransition = 11'd425;
      13: stateTransition = 11'd666;
      14: stateTransition = 11'd425;
      15: stateTransition = 11'd425;
      16: stateTransition = 11'd425;
      17: stateTransition = 11'd425;
      18: stateTransition = 11'd425;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd425;
      22: stateTransition = 11'd425;
      23: stateTransition = 11'd425;
      24: stateTransition = 11'd425;
      25: stateTransition = 11'd425;
      26: stateTransition = 11'd425;
      27: stateTransition = 11'd425;
      28: stateTransition = 11'd425;
      29: stateTransition = 11'd425;
      30: stateTransition = 11'd425;
      31: stateTransition = 11'd425;
      32: stateTransition = 11'd425;
      33: stateTransition = 11'd425;
      34: stateTransition = 11'd425;
      35: stateTransition = 11'd425;
      36: stateTransition = 11'd425;
      37: stateTransition = 11'd425;
      38: stateTransition = 11'd425;
      39: stateTransition = 11'd425;
      40: stateTransition = 11'd425;
      default: stateTransition = 11'bX;
    endcase
    431: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd427;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    432: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd434;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    433: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd447;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    434: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd450;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    435: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd458;
      2: stateTransition = 11'd458;
      3: stateTransition = 11'd458;
      4: stateTransition = 11'd458;
      5: stateTransition = 11'd458;
      6: stateTransition = 11'd458;
      7: stateTransition = 11'd458;
      8: stateTransition = 11'd458;
      9: stateTransition = 11'd432;
      10: stateTransition = 11'd458;
      11: stateTransition = 11'd458;
      12: stateTransition = 11'd458;
      13: stateTransition = 11'd458;
      14: stateTransition = 11'd458;
      15: stateTransition = 11'd458;
      16: stateTransition = 11'd458;
      17: stateTransition = 11'd458;
      18: stateTransition = 11'd458;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd458;
      22: stateTransition = 11'd458;
      23: stateTransition = 11'd458;
      24: stateTransition = 11'd458;
      25: stateTransition = 11'd458;
      26: stateTransition = 11'd458;
      27: stateTransition = 11'd458;
      28: stateTransition = 11'd458;
      29: stateTransition = 11'd458;
      30: stateTransition = 11'd458;
      31: stateTransition = 11'd458;
      32: stateTransition = 11'd458;
      33: stateTransition = 11'd458;
      34: stateTransition = 11'd458;
      35: stateTransition = 11'd458;
      36: stateTransition = 11'd458;
      37: stateTransition = 11'd458;
      38: stateTransition = 11'd458;
      39: stateTransition = 11'd458;
      40: stateTransition = 11'd458;
      default: stateTransition = 11'bX;
    endcase
    436: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd451;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    437: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd446;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    438: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    439: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd425;
      2: stateTransition = 11'd425;
      3: stateTransition = 11'd425;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd437;
      8: stateTransition = 11'd425;
      9: stateTransition = 11'd425;
      10: stateTransition = 11'd425;
      11: stateTransition = 11'd425;
      12: stateTransition = 11'd425;
      13: stateTransition = 11'd666;
      14: stateTransition = 11'd425;
      15: stateTransition = 11'd425;
      16: stateTransition = 11'd425;
      17: stateTransition = 11'd425;
      18: stateTransition = 11'd425;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd440;
      22: stateTransition = 11'd425;
      23: stateTransition = 11'd425;
      24: stateTransition = 11'd442;
      25: stateTransition = 11'd425;
      26: stateTransition = 11'd425;
      27: stateTransition = 11'd425;
      28: stateTransition = 11'd425;
      29: stateTransition = 11'd425;
      30: stateTransition = 11'd425;
      31: stateTransition = 11'd425;
      32: stateTransition = 11'd425;
      33: stateTransition = 11'd425;
      34: stateTransition = 11'd425;
      35: stateTransition = 11'd425;
      36: stateTransition = 11'd425;
      37: stateTransition = 11'd425;
      38: stateTransition = 11'd425;
      39: stateTransition = 11'd425;
      40: stateTransition = 11'd425;
      default: stateTransition = 11'bX;
    endcase
    440: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd438;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    441: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd468;
      2: stateTransition = 11'd468;
      3: stateTransition = 11'd468;
      4: stateTransition = 11'd468;
      5: stateTransition = 11'd468;
      6: stateTransition = 11'd468;
      7: stateTransition = 11'd468;
      8: stateTransition = 11'd468;
      9: stateTransition = 11'd468;
      10: stateTransition = 11'd468;
      11: stateTransition = 11'd468;
      12: stateTransition = 11'd468;
      13: stateTransition = 11'd468;
      14: stateTransition = 11'd468;
      15: stateTransition = 11'd468;
      16: stateTransition = 11'd468;
      17: stateTransition = 11'd468;
      18: stateTransition = 11'd468;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd468;
      22: stateTransition = 11'd468;
      23: stateTransition = 11'd468;
      24: stateTransition = 11'd468;
      25: stateTransition = 11'd468;
      26: stateTransition = 11'd468;
      27: stateTransition = 11'd468;
      28: stateTransition = 11'd468;
      29: stateTransition = 11'd468;
      30: stateTransition = 11'd468;
      31: stateTransition = 11'd468;
      32: stateTransition = 11'd468;
      33: stateTransition = 11'd468;
      34: stateTransition = 11'd468;
      35: stateTransition = 11'd468;
      36: stateTransition = 11'd468;
      37: stateTransition = 11'd468;
      38: stateTransition = 11'd468;
      39: stateTransition = 11'd468;
      40: stateTransition = 11'd468;
      default: stateTransition = 11'bX;
    endcase
    442: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd441;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    443: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd446;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    444: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd454;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    445: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd462;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    446: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd463;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    447: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd458;
      2: stateTransition = 11'd458;
      3: stateTransition = 11'd458;
      4: stateTransition = 11'd458;
      5: stateTransition = 11'd458;
      6: stateTransition = 11'd458;
      7: stateTransition = 11'd458;
      8: stateTransition = 11'd458;
      9: stateTransition = 11'd458;
      10: stateTransition = 11'd458;
      11: stateTransition = 11'd458;
      12: stateTransition = 11'd458;
      13: stateTransition = 11'd458;
      14: stateTransition = 11'd458;
      15: stateTransition = 11'd458;
      16: stateTransition = 11'd458;
      17: stateTransition = 11'd458;
      18: stateTransition = 11'd458;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd458;
      22: stateTransition = 11'd458;
      23: stateTransition = 11'd458;
      24: stateTransition = 11'd458;
      25: stateTransition = 11'd458;
      26: stateTransition = 11'd458;
      27: stateTransition = 11'd458;
      28: stateTransition = 11'd458;
      29: stateTransition = 11'd458;
      30: stateTransition = 11'd458;
      31: stateTransition = 11'd458;
      32: stateTransition = 11'd458;
      33: stateTransition = 11'd458;
      34: stateTransition = 11'd458;
      35: stateTransition = 11'd458;
      36: stateTransition = 11'd458;
      37: stateTransition = 11'd458;
      38: stateTransition = 11'd458;
      39: stateTransition = 11'd458;
      40: stateTransition = 11'd458;
      default: stateTransition = 11'bX;
    endcase
    448: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    449: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd461;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    450: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd457;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    451: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd459;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd480;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    452: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd461;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    453: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd471;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    454: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd467;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    455: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd492;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    456: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd473;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    457: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    458: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd471;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    459: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd469;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    460: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd470;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    461: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd477;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    462: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    463: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd480;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    464: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd189;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd480;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    465: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd502;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    466: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd485;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    467: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd486;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    468: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd487;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    469: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd478;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    470: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd479;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    471: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd480;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    472: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    473: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd492;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    474: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd22;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    475: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd494;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    476: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd495;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    477: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd496;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    478: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd497;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    479: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    480: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd499;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    481: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd501;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    482: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd489;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd609;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    483: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd490;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    484: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd505;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    485: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd504;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    486: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd506;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    487: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd507;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    488: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd508;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    489: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd509;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    490: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd510;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    491: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd511;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    492: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd512;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    493: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd513;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    494: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd514;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    495: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd515;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    496: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd516;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    497: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd517;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    498: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd518;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd686;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    499: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd519;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    500: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd520;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    501: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd521;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    502: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd522;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    503: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd523;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    504: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd523;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    505: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd524;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    506: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd525;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    507: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd528;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    508: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd529;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    509: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd530;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    510: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd526;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    511: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd531;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    512: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd207;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd207;
      9: stateTransition = 11'd533;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd207;
      13: stateTransition = 11'd576;
      14: stateTransition = 11'd207;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd207;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd207;
      22: stateTransition = 11'd207;
      23: stateTransition = 11'd207;
      24: stateTransition = 11'd207;
      25: stateTransition = 11'd207;
      26: stateTransition = 11'd207;
      27: stateTransition = 11'd207;
      28: stateTransition = 11'd207;
      29: stateTransition = 11'd207;
      30: stateTransition = 11'd207;
      31: stateTransition = 11'd207;
      32: stateTransition = 11'd207;
      33: stateTransition = 11'd207;
      34: stateTransition = 11'd207;
      35: stateTransition = 11'd207;
      36: stateTransition = 11'd207;
      37: stateTransition = 11'd207;
      38: stateTransition = 11'd207;
      39: stateTransition = 11'd207;
      40: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    513: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd252;
      2: stateTransition = 11'd252;
      3: stateTransition = 11'd252;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd252;
      8: stateTransition = 11'd534;
      9: stateTransition = 11'd252;
      10: stateTransition = 11'd252;
      11: stateTransition = 11'd252;
      12: stateTransition = 11'd252;
      13: stateTransition = 11'd567;
      14: stateTransition = 11'd252;
      15: stateTransition = 11'd252;
      16: stateTransition = 11'd252;
      17: stateTransition = 11'd252;
      18: stateTransition = 11'd252;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd252;
      22: stateTransition = 11'd252;
      23: stateTransition = 11'd252;
      24: stateTransition = 11'd252;
      25: stateTransition = 11'd252;
      26: stateTransition = 11'd252;
      27: stateTransition = 11'd252;
      28: stateTransition = 11'd252;
      29: stateTransition = 11'd252;
      30: stateTransition = 11'd252;
      31: stateTransition = 11'd252;
      32: stateTransition = 11'd252;
      33: stateTransition = 11'd252;
      34: stateTransition = 11'd252;
      35: stateTransition = 11'd252;
      36: stateTransition = 11'd252;
      37: stateTransition = 11'd252;
      38: stateTransition = 11'd252;
      39: stateTransition = 11'd252;
      40: stateTransition = 11'd252;
      default: stateTransition = 11'bX;
    endcase
    514: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd292;
      2: stateTransition = 11'd535;
      3: stateTransition = 11'd292;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd292;
      8: stateTransition = 11'd292;
      9: stateTransition = 11'd292;
      10: stateTransition = 11'd292;
      11: stateTransition = 11'd292;
      12: stateTransition = 11'd292;
      13: stateTransition = 11'd558;
      14: stateTransition = 11'd292;
      15: stateTransition = 11'd292;
      16: stateTransition = 11'd292;
      17: stateTransition = 11'd292;
      18: stateTransition = 11'd292;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd292;
      22: stateTransition = 11'd292;
      23: stateTransition = 11'd292;
      24: stateTransition = 11'd292;
      25: stateTransition = 11'd292;
      26: stateTransition = 11'd292;
      27: stateTransition = 11'd292;
      28: stateTransition = 11'd292;
      29: stateTransition = 11'd292;
      30: stateTransition = 11'd292;
      31: stateTransition = 11'd292;
      32: stateTransition = 11'd292;
      33: stateTransition = 11'd292;
      34: stateTransition = 11'd292;
      35: stateTransition = 11'd292;
      36: stateTransition = 11'd292;
      37: stateTransition = 11'd292;
      38: stateTransition = 11'd292;
      39: stateTransition = 11'd292;
      40: stateTransition = 11'd292;
      default: stateTransition = 11'bX;
    endcase
    515: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd526;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    516: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd527;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    517: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd329;
      2: stateTransition = 11'd329;
      3: stateTransition = 11'd329;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd329;
      8: stateTransition = 11'd329;
      9: stateTransition = 11'd329;
      10: stateTransition = 11'd329;
      11: stateTransition = 11'd329;
      12: stateTransition = 11'd329;
      13: stateTransition = 11'd548;
      14: stateTransition = 11'd536;
      15: stateTransition = 11'd329;
      16: stateTransition = 11'd329;
      17: stateTransition = 11'd329;
      18: stateTransition = 11'd329;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd329;
      22: stateTransition = 11'd329;
      23: stateTransition = 11'd329;
      24: stateTransition = 11'd329;
      25: stateTransition = 11'd329;
      26: stateTransition = 11'd329;
      27: stateTransition = 11'd329;
      28: stateTransition = 11'd329;
      29: stateTransition = 11'd329;
      30: stateTransition = 11'd329;
      31: stateTransition = 11'd329;
      32: stateTransition = 11'd329;
      33: stateTransition = 11'd329;
      34: stateTransition = 11'd329;
      35: stateTransition = 11'd329;
      36: stateTransition = 11'd329;
      37: stateTransition = 11'd329;
      38: stateTransition = 11'd329;
      39: stateTransition = 11'd329;
      40: stateTransition = 11'd329;
      default: stateTransition = 11'bX;
    endcase
    518: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd532;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    519: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd540;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    520: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd541;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    521: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd542;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    522: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd537;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    523: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd170;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd543;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    524: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd207;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd545;
      9: stateTransition = 11'd207;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd207;
      13: stateTransition = 11'd576;
      14: stateTransition = 11'd207;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd207;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd207;
      22: stateTransition = 11'd207;
      23: stateTransition = 11'd207;
      24: stateTransition = 11'd207;
      25: stateTransition = 11'd207;
      26: stateTransition = 11'd207;
      27: stateTransition = 11'd207;
      28: stateTransition = 11'd207;
      29: stateTransition = 11'd207;
      30: stateTransition = 11'd207;
      31: stateTransition = 11'd207;
      32: stateTransition = 11'd207;
      33: stateTransition = 11'd207;
      34: stateTransition = 11'd207;
      35: stateTransition = 11'd207;
      36: stateTransition = 11'd207;
      37: stateTransition = 11'd207;
      38: stateTransition = 11'd207;
      39: stateTransition = 11'd207;
      40: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    525: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd252;
      2: stateTransition = 11'd546;
      3: stateTransition = 11'd252;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd252;
      8: stateTransition = 11'd252;
      9: stateTransition = 11'd252;
      10: stateTransition = 11'd252;
      11: stateTransition = 11'd252;
      12: stateTransition = 11'd252;
      13: stateTransition = 11'd567;
      14: stateTransition = 11'd252;
      15: stateTransition = 11'd252;
      16: stateTransition = 11'd252;
      17: stateTransition = 11'd252;
      18: stateTransition = 11'd252;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd252;
      22: stateTransition = 11'd252;
      23: stateTransition = 11'd252;
      24: stateTransition = 11'd252;
      25: stateTransition = 11'd252;
      26: stateTransition = 11'd252;
      27: stateTransition = 11'd252;
      28: stateTransition = 11'd252;
      29: stateTransition = 11'd252;
      30: stateTransition = 11'd252;
      31: stateTransition = 11'd252;
      32: stateTransition = 11'd252;
      33: stateTransition = 11'd252;
      34: stateTransition = 11'd252;
      35: stateTransition = 11'd252;
      36: stateTransition = 11'd252;
      37: stateTransition = 11'd252;
      38: stateTransition = 11'd252;
      39: stateTransition = 11'd252;
      40: stateTransition = 11'd252;
      default: stateTransition = 11'bX;
    endcase
    526: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd292;
      2: stateTransition = 11'd292;
      3: stateTransition = 11'd292;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd292;
      8: stateTransition = 11'd292;
      9: stateTransition = 11'd292;
      10: stateTransition = 11'd292;
      11: stateTransition = 11'd292;
      12: stateTransition = 11'd292;
      13: stateTransition = 11'd558;
      14: stateTransition = 11'd547;
      15: stateTransition = 11'd292;
      16: stateTransition = 11'd292;
      17: stateTransition = 11'd292;
      18: stateTransition = 11'd292;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd292;
      22: stateTransition = 11'd292;
      23: stateTransition = 11'd292;
      24: stateTransition = 11'd292;
      25: stateTransition = 11'd292;
      26: stateTransition = 11'd292;
      27: stateTransition = 11'd292;
      28: stateTransition = 11'd292;
      29: stateTransition = 11'd292;
      30: stateTransition = 11'd292;
      31: stateTransition = 11'd292;
      32: stateTransition = 11'd292;
      33: stateTransition = 11'd292;
      34: stateTransition = 11'd292;
      35: stateTransition = 11'd292;
      36: stateTransition = 11'd292;
      37: stateTransition = 11'd292;
      38: stateTransition = 11'd292;
      39: stateTransition = 11'd292;
      40: stateTransition = 11'd292;
      default: stateTransition = 11'bX;
    endcase
    527: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd537;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    528: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd538;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    529: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd544;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    530: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd551;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    531: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd552;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    532: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd553;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    533: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd549;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    534: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd170;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd554;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    535: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd556;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd207;
      9: stateTransition = 11'd207;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd207;
      13: stateTransition = 11'd576;
      14: stateTransition = 11'd207;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd207;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd207;
      22: stateTransition = 11'd207;
      23: stateTransition = 11'd207;
      24: stateTransition = 11'd207;
      25: stateTransition = 11'd207;
      26: stateTransition = 11'd207;
      27: stateTransition = 11'd207;
      28: stateTransition = 11'd207;
      29: stateTransition = 11'd207;
      30: stateTransition = 11'd207;
      31: stateTransition = 11'd207;
      32: stateTransition = 11'd207;
      33: stateTransition = 11'd207;
      34: stateTransition = 11'd207;
      35: stateTransition = 11'd207;
      36: stateTransition = 11'd207;
      37: stateTransition = 11'd207;
      38: stateTransition = 11'd207;
      39: stateTransition = 11'd207;
      40: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    536: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd252;
      2: stateTransition = 11'd252;
      3: stateTransition = 11'd252;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd252;
      8: stateTransition = 11'd252;
      9: stateTransition = 11'd252;
      10: stateTransition = 11'd252;
      11: stateTransition = 11'd252;
      12: stateTransition = 11'd252;
      13: stateTransition = 11'd567;
      14: stateTransition = 11'd557;
      15: stateTransition = 11'd252;
      16: stateTransition = 11'd252;
      17: stateTransition = 11'd252;
      18: stateTransition = 11'd252;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd252;
      22: stateTransition = 11'd252;
      23: stateTransition = 11'd252;
      24: stateTransition = 11'd252;
      25: stateTransition = 11'd252;
      26: stateTransition = 11'd252;
      27: stateTransition = 11'd252;
      28: stateTransition = 11'd252;
      29: stateTransition = 11'd252;
      30: stateTransition = 11'd252;
      31: stateTransition = 11'd252;
      32: stateTransition = 11'd252;
      33: stateTransition = 11'd252;
      34: stateTransition = 11'd252;
      35: stateTransition = 11'd252;
      36: stateTransition = 11'd252;
      37: stateTransition = 11'd252;
      38: stateTransition = 11'd252;
      39: stateTransition = 11'd252;
      40: stateTransition = 11'd252;
      default: stateTransition = 11'bX;
    endcase
    537: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd549;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    538: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd550;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    539: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd555;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    540: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd561;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    541: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd562;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    542: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd563;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    543: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd559;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    544: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd564;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd170;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    545: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd207;
      2: stateTransition = 11'd207;
      3: stateTransition = 11'd207;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd207;
      8: stateTransition = 11'd207;
      9: stateTransition = 11'd207;
      10: stateTransition = 11'd207;
      11: stateTransition = 11'd207;
      12: stateTransition = 11'd207;
      13: stateTransition = 11'd576;
      14: stateTransition = 11'd566;
      15: stateTransition = 11'd207;
      16: stateTransition = 11'd207;
      17: stateTransition = 11'd207;
      18: stateTransition = 11'd207;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd207;
      22: stateTransition = 11'd207;
      23: stateTransition = 11'd207;
      24: stateTransition = 11'd207;
      25: stateTransition = 11'd207;
      26: stateTransition = 11'd207;
      27: stateTransition = 11'd207;
      28: stateTransition = 11'd207;
      29: stateTransition = 11'd207;
      30: stateTransition = 11'd207;
      31: stateTransition = 11'd207;
      32: stateTransition = 11'd207;
      33: stateTransition = 11'd207;
      34: stateTransition = 11'd207;
      35: stateTransition = 11'd207;
      36: stateTransition = 11'd207;
      37: stateTransition = 11'd207;
      38: stateTransition = 11'd207;
      39: stateTransition = 11'd207;
      40: stateTransition = 11'd207;
      default: stateTransition = 11'bX;
    endcase
    546: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd560;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    547: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd559;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    548: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd560;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    549: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd565;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    550: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd571;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    551: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd572;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    552: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd573;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd126;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    553: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd569;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    554: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd170;
      2: stateTransition = 11'd170;
      3: stateTransition = 11'd170;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd170;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd170;
      10: stateTransition = 11'd170;
      11: stateTransition = 11'd170;
      12: stateTransition = 11'd170;
      13: stateTransition = 11'd584;
      14: stateTransition = 11'd574;
      15: stateTransition = 11'd170;
      16: stateTransition = 11'd170;
      17: stateTransition = 11'd170;
      18: stateTransition = 11'd170;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd170;
      22: stateTransition = 11'd170;
      23: stateTransition = 11'd170;
      24: stateTransition = 11'd170;
      25: stateTransition = 11'd170;
      26: stateTransition = 11'd170;
      27: stateTransition = 11'd170;
      28: stateTransition = 11'd170;
      29: stateTransition = 11'd170;
      30: stateTransition = 11'd170;
      31: stateTransition = 11'd170;
      32: stateTransition = 11'd170;
      33: stateTransition = 11'd170;
      34: stateTransition = 11'd170;
      35: stateTransition = 11'd170;
      36: stateTransition = 11'd170;
      37: stateTransition = 11'd170;
      38: stateTransition = 11'd170;
      39: stateTransition = 11'd170;
      40: stateTransition = 11'd170;
      default: stateTransition = 11'bX;
    endcase
    555: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd568;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    556: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd570;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    557: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd569;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    558: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd570;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    559: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd575;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    560: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd581;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    561: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd582;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd64;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    562: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd126;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd126;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd126;
      9: stateTransition = 11'd126;
      10: stateTransition = 11'd126;
      11: stateTransition = 11'd126;
      12: stateTransition = 11'd126;
      13: stateTransition = 11'd593;
      14: stateTransition = 11'd583;
      15: stateTransition = 11'd126;
      16: stateTransition = 11'd126;
      17: stateTransition = 11'd126;
      18: stateTransition = 11'd126;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd126;
      22: stateTransition = 11'd126;
      23: stateTransition = 11'd126;
      24: stateTransition = 11'd126;
      25: stateTransition = 11'd126;
      26: stateTransition = 11'd126;
      27: stateTransition = 11'd126;
      28: stateTransition = 11'd126;
      29: stateTransition = 11'd126;
      30: stateTransition = 11'd126;
      31: stateTransition = 11'd126;
      32: stateTransition = 11'd126;
      33: stateTransition = 11'd126;
      34: stateTransition = 11'd126;
      35: stateTransition = 11'd126;
      36: stateTransition = 11'd126;
      37: stateTransition = 11'd126;
      38: stateTransition = 11'd126;
      39: stateTransition = 11'd126;
      40: stateTransition = 11'd126;
      default: stateTransition = 11'bX;
    endcase
    563: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd579;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    564: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd577;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    565: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd578;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    566: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd580;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    567: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd579;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    568: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd580;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    569: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd585;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    570: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd591;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd24;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    571: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd64;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd64;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd64;
      8: stateTransition = 11'd64;
      9: stateTransition = 11'd64;
      10: stateTransition = 11'd64;
      11: stateTransition = 11'd64;
      12: stateTransition = 11'd64;
      13: stateTransition = 11'd602;
      14: stateTransition = 11'd592;
      15: stateTransition = 11'd64;
      16: stateTransition = 11'd64;
      17: stateTransition = 11'd64;
      18: stateTransition = 11'd64;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd64;
      22: stateTransition = 11'd64;
      23: stateTransition = 11'd64;
      24: stateTransition = 11'd64;
      25: stateTransition = 11'd64;
      26: stateTransition = 11'd64;
      27: stateTransition = 11'd64;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd64;
      30: stateTransition = 11'd64;
      31: stateTransition = 11'd64;
      32: stateTransition = 11'd64;
      33: stateTransition = 11'd64;
      34: stateTransition = 11'd64;
      35: stateTransition = 11'd64;
      36: stateTransition = 11'd64;
      37: stateTransition = 11'd64;
      38: stateTransition = 11'd64;
      39: stateTransition = 11'd64;
      40: stateTransition = 11'd64;
      default: stateTransition = 11'bX;
    endcase
    572: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd589;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    573: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd586;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    574: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd587;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    575: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd588;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    576: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd590;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    577: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd589;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    578: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd590;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    579: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd594;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd172;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    580: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd24;
      2: stateTransition = 11'd24;
      3: stateTransition = 11'd24;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd24;
      8: stateTransition = 11'd24;
      9: stateTransition = 11'd24;
      10: stateTransition = 11'd24;
      11: stateTransition = 11'd24;
      12: stateTransition = 11'd24;
      13: stateTransition = 11'd611;
      14: stateTransition = 11'd601;
      15: stateTransition = 11'd24;
      16: stateTransition = 11'd24;
      17: stateTransition = 11'd24;
      18: stateTransition = 11'd24;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd24;
      22: stateTransition = 11'd24;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd24;
      25: stateTransition = 11'd24;
      26: stateTransition = 11'd24;
      27: stateTransition = 11'd24;
      28: stateTransition = 11'd24;
      29: stateTransition = 11'd24;
      30: stateTransition = 11'd24;
      31: stateTransition = 11'd24;
      32: stateTransition = 11'd24;
      33: stateTransition = 11'd24;
      34: stateTransition = 11'd24;
      35: stateTransition = 11'd24;
      36: stateTransition = 11'd24;
      37: stateTransition = 11'd24;
      38: stateTransition = 11'd24;
      39: stateTransition = 11'd24;
      40: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    581: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd599;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    582: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd595;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    583: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd596;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    584: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd597;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    585: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd598;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    586: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd600;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    587: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd599;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd503;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    588: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd600;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    589: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd172;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd172;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd172;
      8: stateTransition = 11'd172;
      9: stateTransition = 11'd172;
      10: stateTransition = 11'd172;
      11: stateTransition = 11'd172;
      12: stateTransition = 11'd172;
      13: stateTransition = 11'd612;
      14: stateTransition = 11'd603;
      15: stateTransition = 11'd172;
      16: stateTransition = 11'd172;
      17: stateTransition = 11'd172;
      18: stateTransition = 11'd172;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd172;
      22: stateTransition = 11'd172;
      23: stateTransition = 11'd172;
      24: stateTransition = 11'd172;
      25: stateTransition = 11'd172;
      26: stateTransition = 11'd172;
      27: stateTransition = 11'd172;
      28: stateTransition = 11'd172;
      29: stateTransition = 11'd172;
      30: stateTransition = 11'd172;
      31: stateTransition = 11'd172;
      32: stateTransition = 11'd172;
      33: stateTransition = 11'd172;
      34: stateTransition = 11'd172;
      35: stateTransition = 11'd172;
      36: stateTransition = 11'd172;
      37: stateTransition = 11'd172;
      38: stateTransition = 11'd172;
      39: stateTransition = 11'd172;
      40: stateTransition = 11'd172;
      default: stateTransition = 11'bX;
    endcase
    590: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd129;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd609;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    591: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd604;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    592: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd605;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    593: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd606;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    594: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd607;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    595: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd608;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    596: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd610;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    597: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd503;
      2: stateTransition = 11'd503;
      3: stateTransition = 11'd503;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd503;
      8: stateTransition = 11'd503;
      9: stateTransition = 11'd503;
      10: stateTransition = 11'd503;
      11: stateTransition = 11'd503;
      12: stateTransition = 11'd503;
      13: stateTransition = 11'd619;
      14: stateTransition = 11'd609;
      15: stateTransition = 11'd503;
      16: stateTransition = 11'd503;
      17: stateTransition = 11'd503;
      18: stateTransition = 11'd503;
      19: stateTransition = 11'd503;
      20: stateTransition = 11'd503;
      21: stateTransition = 11'd503;
      22: stateTransition = 11'd503;
      23: stateTransition = 11'd503;
      24: stateTransition = 11'd503;
      25: stateTransition = 11'd503;
      26: stateTransition = 11'd503;
      27: stateTransition = 11'd503;
      28: stateTransition = 11'd503;
      29: stateTransition = 11'd503;
      30: stateTransition = 11'd503;
      31: stateTransition = 11'd503;
      32: stateTransition = 11'd503;
      33: stateTransition = 11'd503;
      34: stateTransition = 11'd503;
      35: stateTransition = 11'd503;
      36: stateTransition = 11'd503;
      37: stateTransition = 11'd503;
      38: stateTransition = 11'd503;
      39: stateTransition = 11'd503;
      40: stateTransition = 11'd503;
      default: stateTransition = 11'bX;
    endcase
    598: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd610;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    599: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd613;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    600: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd614;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    601: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd615;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    602: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd616;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    603: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd617;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    604: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd618;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    605: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd620;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    606: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd620;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    607: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd621;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    608: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd622;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    609: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd623;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    610: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd624;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    611: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd625;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    612: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd626;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    613: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd627;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    614: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd628;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    615: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd628;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    616: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd629;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    617: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd630;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    618: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd631;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    619: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd632;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    620: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd633;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    621: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd634;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    622: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd635;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    623: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd636;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    624: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd637;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    625: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd637;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    626: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd638;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    627: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd639;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    628: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd648;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    629: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd640;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    630: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd650;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd677;
      14: stateTransition = 11'd399;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd399;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd399;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd399;
      35: stateTransition = 11'd399;
      36: stateTransition = 11'd399;
      37: stateTransition = 11'd399;
      38: stateTransition = 11'd399;
      39: stateTransition = 11'd399;
      40: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    631: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd641;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    632: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd425;
      2: stateTransition = 11'd425;
      3: stateTransition = 11'd425;
      4: stateTransition = 11'd460;
      5: stateTransition = 11'd460;
      6: stateTransition = 11'd460;
      7: stateTransition = 11'd437;
      8: stateTransition = 11'd425;
      9: stateTransition = 11'd425;
      10: stateTransition = 11'd425;
      11: stateTransition = 11'd425;
      12: stateTransition = 11'd425;
      13: stateTransition = 11'd666;
      14: stateTransition = 11'd652;
      15: stateTransition = 11'd425;
      16: stateTransition = 11'd425;
      17: stateTransition = 11'd425;
      18: stateTransition = 11'd425;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd425;
      22: stateTransition = 11'd425;
      23: stateTransition = 11'd425;
      24: stateTransition = 11'd425;
      25: stateTransition = 11'd425;
      26: stateTransition = 11'd425;
      27: stateTransition = 11'd425;
      28: stateTransition = 11'd425;
      29: stateTransition = 11'd425;
      30: stateTransition = 11'd425;
      31: stateTransition = 11'd425;
      32: stateTransition = 11'd425;
      33: stateTransition = 11'd425;
      34: stateTransition = 11'd425;
      35: stateTransition = 11'd425;
      36: stateTransition = 11'd425;
      37: stateTransition = 11'd425;
      38: stateTransition = 11'd425;
      39: stateTransition = 11'd425;
      40: stateTransition = 11'd425;
      default: stateTransition = 11'bX;
    endcase
    633: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd642;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    634: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd643;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    635: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd644;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    636: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd645;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    637: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd646;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    638: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd647;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    639: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd647;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    640: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd649;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    641: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd651;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    642: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd662;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd369;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    643: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd653;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    644: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd399;
      2: stateTransition = 11'd399;
      3: stateTransition = 11'd399;
      4: stateTransition = 11'd439;
      5: stateTransition = 11'd439;
      6: stateTransition = 11'd439;
      7: stateTransition = 11'd413;
      8: stateTransition = 11'd399;
      9: stateTransition = 11'd399;
      10: stateTransition = 11'd399;
      11: stateTransition = 11'd399;
      12: stateTransition = 11'd399;
      13: stateTransition = 11'd677;
      14: stateTransition = 11'd664;
      15: stateTransition = 11'd399;
      16: stateTransition = 11'd399;
      17: stateTransition = 11'd399;
      18: stateTransition = 11'd399;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd399;
      22: stateTransition = 11'd399;
      23: stateTransition = 11'd399;
      24: stateTransition = 11'd399;
      25: stateTransition = 11'd399;
      26: stateTransition = 11'd399;
      27: stateTransition = 11'd399;
      28: stateTransition = 11'd399;
      29: stateTransition = 11'd399;
      30: stateTransition = 11'd399;
      31: stateTransition = 11'd399;
      32: stateTransition = 11'd399;
      33: stateTransition = 11'd399;
      34: stateTransition = 11'd399;
      35: stateTransition = 11'd399;
      36: stateTransition = 11'd399;
      37: stateTransition = 11'd399;
      38: stateTransition = 11'd399;
      39: stateTransition = 11'd399;
      40: stateTransition = 11'd399;
      default: stateTransition = 11'bX;
    endcase
    645: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd655;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    646: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd656;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    647: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd657;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    648: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd658;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    649: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd659;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    650: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd660;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    651: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd661;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    652: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd661;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    653: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd663;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd383;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    654: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd665;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd411;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    655: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd369;
      2: stateTransition = 11'd369;
      3: stateTransition = 11'd369;
      4: stateTransition = 11'd421;
      5: stateTransition = 11'd421;
      6: stateTransition = 11'd421;
      7: stateTransition = 11'd385;
      8: stateTransition = 11'd369;
      9: stateTransition = 11'd369;
      10: stateTransition = 11'd369;
      11: stateTransition = 11'd369;
      12: stateTransition = 11'd369;
      13: stateTransition = 11'd688;
      14: stateTransition = 11'd675;
      15: stateTransition = 11'd369;
      16: stateTransition = 11'd369;
      17: stateTransition = 11'd369;
      18: stateTransition = 11'd369;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd369;
      22: stateTransition = 11'd369;
      23: stateTransition = 11'd369;
      24: stateTransition = 11'd369;
      25: stateTransition = 11'd369;
      26: stateTransition = 11'd369;
      27: stateTransition = 11'd369;
      28: stateTransition = 11'd369;
      29: stateTransition = 11'd369;
      30: stateTransition = 11'd369;
      31: stateTransition = 11'd369;
      32: stateTransition = 11'd369;
      33: stateTransition = 11'd369;
      34: stateTransition = 11'd369;
      35: stateTransition = 11'd369;
      36: stateTransition = 11'd369;
      37: stateTransition = 11'd369;
      38: stateTransition = 11'd369;
      39: stateTransition = 11'd369;
      40: stateTransition = 11'd369;
      default: stateTransition = 11'bX;
    endcase
    656: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd667;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd436;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    657: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd668;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd455;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    658: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd669;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd466;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    659: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd670;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd476;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    660: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd671;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd482;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    661: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd672;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd493;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    662: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd673;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd500;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    663: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd674;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    664: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd674;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd13;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    665: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd189;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd686;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    666: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd383;
      2: stateTransition = 11'd383;
      3: stateTransition = 11'd383;
      4: stateTransition = 11'd393;
      5: stateTransition = 11'd393;
      6: stateTransition = 11'd393;
      7: stateTransition = 11'd353;
      8: stateTransition = 11'd383;
      9: stateTransition = 11'd383;
      10: stateTransition = 11'd383;
      11: stateTransition = 11'd383;
      12: stateTransition = 11'd383;
      13: stateTransition = 11'd689;
      14: stateTransition = 11'd676;
      15: stateTransition = 11'd383;
      16: stateTransition = 11'd383;
      17: stateTransition = 11'd383;
      18: stateTransition = 11'd383;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd383;
      22: stateTransition = 11'd383;
      23: stateTransition = 11'd383;
      24: stateTransition = 11'd383;
      25: stateTransition = 11'd383;
      26: stateTransition = 11'd383;
      27: stateTransition = 11'd383;
      28: stateTransition = 11'd383;
      29: stateTransition = 11'd383;
      30: stateTransition = 11'd383;
      31: stateTransition = 11'd383;
      32: stateTransition = 11'd383;
      33: stateTransition = 11'd383;
      34: stateTransition = 11'd383;
      35: stateTransition = 11'd383;
      36: stateTransition = 11'd383;
      37: stateTransition = 11'd383;
      38: stateTransition = 11'd383;
      39: stateTransition = 11'd383;
      40: stateTransition = 11'd383;
      default: stateTransition = 11'bX;
    endcase
    667: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd411;
      2: stateTransition = 11'd411;
      3: stateTransition = 11'd411;
      4: stateTransition = 11'd358;
      5: stateTransition = 11'd358;
      6: stateTransition = 11'd358;
      7: stateTransition = 11'd382;
      8: stateTransition = 11'd411;
      9: stateTransition = 11'd411;
      10: stateTransition = 11'd411;
      11: stateTransition = 11'd411;
      12: stateTransition = 11'd411;
      13: stateTransition = 11'd690;
      14: stateTransition = 11'd678;
      15: stateTransition = 11'd411;
      16: stateTransition = 11'd411;
      17: stateTransition = 11'd411;
      18: stateTransition = 11'd411;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd411;
      22: stateTransition = 11'd411;
      23: stateTransition = 11'd411;
      24: stateTransition = 11'd411;
      25: stateTransition = 11'd411;
      26: stateTransition = 11'd411;
      27: stateTransition = 11'd411;
      28: stateTransition = 11'd411;
      29: stateTransition = 11'd411;
      30: stateTransition = 11'd411;
      31: stateTransition = 11'd411;
      32: stateTransition = 11'd411;
      33: stateTransition = 11'd411;
      34: stateTransition = 11'd411;
      35: stateTransition = 11'd411;
      36: stateTransition = 11'd411;
      37: stateTransition = 11'd411;
      38: stateTransition = 11'd411;
      39: stateTransition = 11'd411;
      40: stateTransition = 11'd411;
      default: stateTransition = 11'bX;
    endcase
    668: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd436;
      2: stateTransition = 11'd436;
      3: stateTransition = 11'd436;
      4: stateTransition = 11'd316;
      5: stateTransition = 11'd316;
      6: stateTransition = 11'd316;
      7: stateTransition = 11'd410;
      8: stateTransition = 11'd436;
      9: stateTransition = 11'd436;
      10: stateTransition = 11'd436;
      11: stateTransition = 11'd436;
      12: stateTransition = 11'd436;
      13: stateTransition = 11'd691;
      14: stateTransition = 11'd679;
      15: stateTransition = 11'd436;
      16: stateTransition = 11'd436;
      17: stateTransition = 11'd436;
      18: stateTransition = 11'd436;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd436;
      22: stateTransition = 11'd436;
      23: stateTransition = 11'd436;
      24: stateTransition = 11'd436;
      25: stateTransition = 11'd436;
      26: stateTransition = 11'd436;
      27: stateTransition = 11'd436;
      28: stateTransition = 11'd436;
      29: stateTransition = 11'd436;
      30: stateTransition = 11'd436;
      31: stateTransition = 11'd436;
      32: stateTransition = 11'd436;
      33: stateTransition = 11'd436;
      34: stateTransition = 11'd436;
      35: stateTransition = 11'd436;
      36: stateTransition = 11'd436;
      37: stateTransition = 11'd436;
      38: stateTransition = 11'd436;
      39: stateTransition = 11'd436;
      40: stateTransition = 11'd436;
      default: stateTransition = 11'bX;
    endcase
    669: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd455;
      2: stateTransition = 11'd455;
      3: stateTransition = 11'd455;
      4: stateTransition = 11'd274;
      5: stateTransition = 11'd274;
      6: stateTransition = 11'd274;
      7: stateTransition = 11'd435;
      8: stateTransition = 11'd455;
      9: stateTransition = 11'd455;
      10: stateTransition = 11'd455;
      11: stateTransition = 11'd455;
      12: stateTransition = 11'd455;
      13: stateTransition = 11'd692;
      14: stateTransition = 11'd680;
      15: stateTransition = 11'd455;
      16: stateTransition = 11'd455;
      17: stateTransition = 11'd455;
      18: stateTransition = 11'd455;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd455;
      22: stateTransition = 11'd455;
      23: stateTransition = 11'd455;
      24: stateTransition = 11'd455;
      25: stateTransition = 11'd455;
      26: stateTransition = 11'd455;
      27: stateTransition = 11'd455;
      28: stateTransition = 11'd455;
      29: stateTransition = 11'd455;
      30: stateTransition = 11'd455;
      31: stateTransition = 11'd455;
      32: stateTransition = 11'd455;
      33: stateTransition = 11'd455;
      34: stateTransition = 11'd455;
      35: stateTransition = 11'd455;
      36: stateTransition = 11'd455;
      37: stateTransition = 11'd455;
      38: stateTransition = 11'd455;
      39: stateTransition = 11'd455;
      40: stateTransition = 11'd455;
      default: stateTransition = 11'bX;
    endcase
    670: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd466;
      2: stateTransition = 11'd466;
      3: stateTransition = 11'd466;
      4: stateTransition = 11'd238;
      5: stateTransition = 11'd238;
      6: stateTransition = 11'd238;
      7: stateTransition = 11'd453;
      8: stateTransition = 11'd466;
      9: stateTransition = 11'd466;
      10: stateTransition = 11'd466;
      11: stateTransition = 11'd466;
      12: stateTransition = 11'd466;
      13: stateTransition = 11'd693;
      14: stateTransition = 11'd681;
      15: stateTransition = 11'd466;
      16: stateTransition = 11'd466;
      17: stateTransition = 11'd466;
      18: stateTransition = 11'd466;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd466;
      22: stateTransition = 11'd466;
      23: stateTransition = 11'd466;
      24: stateTransition = 11'd466;
      25: stateTransition = 11'd466;
      26: stateTransition = 11'd466;
      27: stateTransition = 11'd466;
      28: stateTransition = 11'd466;
      29: stateTransition = 11'd466;
      30: stateTransition = 11'd466;
      31: stateTransition = 11'd466;
      32: stateTransition = 11'd466;
      33: stateTransition = 11'd466;
      34: stateTransition = 11'd466;
      35: stateTransition = 11'd466;
      36: stateTransition = 11'd466;
      37: stateTransition = 11'd466;
      38: stateTransition = 11'd466;
      39: stateTransition = 11'd466;
      40: stateTransition = 11'd466;
      default: stateTransition = 11'bX;
    endcase
    671: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd476;
      2: stateTransition = 11'd476;
      3: stateTransition = 11'd476;
      4: stateTransition = 11'd186;
      5: stateTransition = 11'd186;
      6: stateTransition = 11'd186;
      7: stateTransition = 11'd464;
      8: stateTransition = 11'd476;
      9: stateTransition = 11'd476;
      10: stateTransition = 11'd476;
      11: stateTransition = 11'd476;
      12: stateTransition = 11'd476;
      13: stateTransition = 11'd694;
      14: stateTransition = 11'd682;
      15: stateTransition = 11'd476;
      16: stateTransition = 11'd476;
      17: stateTransition = 11'd476;
      18: stateTransition = 11'd476;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd476;
      22: stateTransition = 11'd476;
      23: stateTransition = 11'd476;
      24: stateTransition = 11'd476;
      25: stateTransition = 11'd476;
      26: stateTransition = 11'd476;
      27: stateTransition = 11'd476;
      28: stateTransition = 11'd476;
      29: stateTransition = 11'd476;
      30: stateTransition = 11'd476;
      31: stateTransition = 11'd476;
      32: stateTransition = 11'd476;
      33: stateTransition = 11'd476;
      34: stateTransition = 11'd476;
      35: stateTransition = 11'd476;
      36: stateTransition = 11'd476;
      37: stateTransition = 11'd476;
      38: stateTransition = 11'd476;
      39: stateTransition = 11'd476;
      40: stateTransition = 11'd476;
      default: stateTransition = 11'bX;
    endcase
    672: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd482;
      2: stateTransition = 11'd482;
      3: stateTransition = 11'd482;
      4: stateTransition = 11'd152;
      5: stateTransition = 11'd152;
      6: stateTransition = 11'd152;
      7: stateTransition = 11'd475;
      8: stateTransition = 11'd482;
      9: stateTransition = 11'd482;
      10: stateTransition = 11'd482;
      11: stateTransition = 11'd482;
      12: stateTransition = 11'd482;
      13: stateTransition = 11'd695;
      14: stateTransition = 11'd683;
      15: stateTransition = 11'd482;
      16: stateTransition = 11'd482;
      17: stateTransition = 11'd482;
      18: stateTransition = 11'd482;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd482;
      22: stateTransition = 11'd482;
      23: stateTransition = 11'd482;
      24: stateTransition = 11'd482;
      25: stateTransition = 11'd482;
      26: stateTransition = 11'd482;
      27: stateTransition = 11'd482;
      28: stateTransition = 11'd482;
      29: stateTransition = 11'd482;
      30: stateTransition = 11'd482;
      31: stateTransition = 11'd482;
      32: stateTransition = 11'd482;
      33: stateTransition = 11'd482;
      34: stateTransition = 11'd482;
      35: stateTransition = 11'd482;
      36: stateTransition = 11'd482;
      37: stateTransition = 11'd482;
      38: stateTransition = 11'd482;
      39: stateTransition = 11'd482;
      40: stateTransition = 11'd482;
      default: stateTransition = 11'bX;
    endcase
    673: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd493;
      2: stateTransition = 11'd493;
      3: stateTransition = 11'd493;
      4: stateTransition = 11'd105;
      5: stateTransition = 11'd105;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd481;
      8: stateTransition = 11'd493;
      9: stateTransition = 11'd493;
      10: stateTransition = 11'd493;
      11: stateTransition = 11'd493;
      12: stateTransition = 11'd493;
      13: stateTransition = 11'd696;
      14: stateTransition = 11'd684;
      15: stateTransition = 11'd493;
      16: stateTransition = 11'd493;
      17: stateTransition = 11'd493;
      18: stateTransition = 11'd493;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd493;
      22: stateTransition = 11'd493;
      23: stateTransition = 11'd493;
      24: stateTransition = 11'd493;
      25: stateTransition = 11'd493;
      26: stateTransition = 11'd493;
      27: stateTransition = 11'd493;
      28: stateTransition = 11'd493;
      29: stateTransition = 11'd493;
      30: stateTransition = 11'd493;
      31: stateTransition = 11'd493;
      32: stateTransition = 11'd493;
      33: stateTransition = 11'd493;
      34: stateTransition = 11'd493;
      35: stateTransition = 11'd493;
      36: stateTransition = 11'd493;
      37: stateTransition = 11'd493;
      38: stateTransition = 11'd493;
      39: stateTransition = 11'd493;
      40: stateTransition = 11'd493;
      default: stateTransition = 11'bX;
    endcase
    674: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd500;
      2: stateTransition = 11'd500;
      3: stateTransition = 11'd500;
      4: stateTransition = 11'd27;
      5: stateTransition = 11'd27;
      6: stateTransition = 11'd27;
      7: stateTransition = 11'd483;
      8: stateTransition = 11'd500;
      9: stateTransition = 11'd500;
      10: stateTransition = 11'd500;
      11: stateTransition = 11'd500;
      12: stateTransition = 11'd500;
      13: stateTransition = 11'd697;
      14: stateTransition = 11'd685;
      15: stateTransition = 11'd500;
      16: stateTransition = 11'd500;
      17: stateTransition = 11'd500;
      18: stateTransition = 11'd500;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd500;
      22: stateTransition = 11'd500;
      23: stateTransition = 11'd500;
      24: stateTransition = 11'd500;
      25: stateTransition = 11'd500;
      26: stateTransition = 11'd500;
      27: stateTransition = 11'd500;
      28: stateTransition = 11'd500;
      29: stateTransition = 11'd500;
      30: stateTransition = 11'd500;
      31: stateTransition = 11'd500;
      32: stateTransition = 11'd500;
      33: stateTransition = 11'd500;
      34: stateTransition = 11'd500;
      35: stateTransition = 11'd500;
      36: stateTransition = 11'd500;
      37: stateTransition = 11'd500;
      38: stateTransition = 11'd500;
      39: stateTransition = 11'd500;
      40: stateTransition = 11'd500;
      default: stateTransition = 11'bX;
    endcase
    675: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd498;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd686;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    676: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd13;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd13;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd491;
      8: stateTransition = 11'd13;
      9: stateTransition = 11'd13;
      10: stateTransition = 11'd13;
      11: stateTransition = 11'd13;
      12: stateTransition = 11'd13;
      13: stateTransition = 11'd698;
      14: stateTransition = 11'd686;
      15: stateTransition = 11'd13;
      16: stateTransition = 11'd13;
      17: stateTransition = 11'd13;
      18: stateTransition = 11'd13;
      19: stateTransition = 11'd13;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd13;
      23: stateTransition = 11'd13;
      24: stateTransition = 11'd13;
      25: stateTransition = 11'd13;
      26: stateTransition = 11'd13;
      27: stateTransition = 11'd13;
      28: stateTransition = 11'd13;
      29: stateTransition = 11'd13;
      30: stateTransition = 11'd13;
      31: stateTransition = 11'd13;
      32: stateTransition = 11'd13;
      33: stateTransition = 11'd13;
      34: stateTransition = 11'd13;
      35: stateTransition = 11'd13;
      36: stateTransition = 11'd13;
      37: stateTransition = 11'd13;
      38: stateTransition = 11'd13;
      39: stateTransition = 11'd13;
      40: stateTransition = 11'd13;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
