   parameter w_din = 32 ,
	       size = 8 ,
	       log2size = 3;
   
