/* ----------------------------------------------------------
 Generalized Descriptor Unpacker (version1: max(field_width) < input data width
 ==========================================================
 Full parameterized:
 
 Parameters: N = width of input bus
             M = width multiplier, output bus width = N*M
             LOG2M = ceiling( log2(M) )
             default: 8 bit ==> 32 bit ,N=8,M=4,LOG2M=2
 
 Examples: 
 
 For self test , compile this file with +define+TEST

 inputs:
   clk   => posedge triggered
   reset => active high
   din   => input data bus
   valid_din => active high, signals valid data on input bus
  
 outputs:
  
 Author: VJ Sananda

---------------------------------------------------------- */

`include "gdu.vh"

module gdu (/*AUTOARG*/
   // Outputs
   err, valid_f0, valid_f1, valid_f2, valid_f3, valid_f4, dout_f0, 
   dout_f1, dout_f2, dout_f3, dout_f4, 
   // Inputs
   clk, reset, sop, eop, din, valid_din
   );

   parameter W = 32 ;//Width of data input bus
   parameter N = 3 ;//Number of data words in packet
   parameter LOG2N = 2 ;//Ceiling of Log2(N)
   
   parameter BIGENDIAN = 0;//1 if big endian
   
   input clk ;
   input reset ;
   input sop ;
   input eop ;

   
   input [W-1:0]   din ;
   input 	   valid_din ;

   output 	   err ;

   // Should be autogenerated based on packet defn
   output valid_f0 ;
   output valid_f1 ;
   output valid_f2 ;
   output valid_f3 ;
   output valid_f4 ;

   output [`F0_W-1:0] dout_f0 ;
   output [`F1_W-1:0] dout_f1 ;
   output [`F2_W-1:0] dout_f2 ;
   output [`F3_W-1:0] dout_f3 ;
   output [`F4_W-1:0] dout_f4 ;

   reg valid_f0 ;
   reg valid_f1 ;
   reg valid_f2 ;
   reg valid_f3 ;
   reg valid_f4 ;

   reg [`F0_W-1:0] dout_f0 ;
   reg [`F1_W-1:0] dout_f1 ;
   reg [`F2_W-1:0] dout_f2 ;
   reg [`F3_W-1:0] dout_f3 ;
   reg [`F4_W-1:0] dout_f4 ;   

   // ---------- END INPUT/OUTPUT DECL ----------

   //---------------------------------------------
   //A note about the suffixes
   //
   //   _[r,w].[c,d].[#] : choose 1 of the letters in each [] and
   //                      concatenate to build suffix
   //
   //[r,w]: r=>register, w=>wire
   //
   //[c,d]: c=>control,  d=>datapath
   //
   //[#] : Number, reflects register stage number
   //Within a clocked always block, signal on the LHS
   //of a non-blocking assignment, will have this number incremented
   //beyond the largest # of the expression on the RHS or that in a
   //conditional expression controlling the assignment
   //
   //On a wire assign, this number will not increment.
   //Goal is to make the clock cycle dependencies obvious
   //---------------------------------------------

   wire [LOG2N-1:0]  cnt_wc1;   
   reg  [LOG2N-1:0]  cnt_rc2;

   reg [W-1:0]	   hold_rd1 ;

   wire 	   end_of_count_wc2 = (cnt_rc2 == N-1);
   
   //Control Counter
   always @(posedge clk or posedge reset)
     //if N is not a power of 2, addcondition to reset
     if (reset || eop || (end_of_count_wc2 & valid_din  )  )
       cnt_rc2 <= 0;
     else
       if ( valid_din )
	 cnt_rc2 <= cnt_wc1;
   assign 	     cnt_wc1 = cnt_rc2 + 1 ;
   
   always @(posedge clk or posedge reset)
     if ( reset )
       begin
	  valid_f0 <= 0;
	  valid_f1 <= 0;
	  valid_f2 <= 0;
	  valid_f3 <= 0;
	  valid_f4 <= 0;	  	  	  
       end
     else
       begin
	  //This section has to be autogenerated from pkt defn
	  valid_f0 <= 0;
	  valid_f1 <= 0;
	  valid_f2 <= 0;
	  valid_f3 <= 0;
	  valid_f4 <= 0;	  	  
	
	  if ( valid_din )
	    begin
	       hold_rd1 <= din ;
	       
	       case(cnt_rc2)
		 0: begin
		    valid_f0 <= 1 ;
		    dout_f0  <= din[`f0_W0_MSB:`f0_W0_LSB] ;
		    valid_f1 <= 1;
		    dout_f1  <= din[`f1_W0_MSB:`f1_W0_LSB];
		 end
		 1: begin
		    valid_f2 <= 1 ;
		    dout_f2  <= { din[`f2_W1_MSB:`f2_W1_LSB] , hold_rd1[`f2_W0_MSB:`f2_W0_LSB] };
		 end
		 2: begin
		    valid_f3 <= 1 ;
		    dout_f3  <= { din[`f3_W2_MSB:`f3_W2_LSB] , hold_rd1[`f3_W1_MSB:`f3_W1_LSB] };
		    valid_f4 <= 1 ;
		    dout_f4  <= din[`f4_W2_MSB:`f4_W2_LSB ];
		 end	 
	       endcase // caseendcase
	    end // if ( valid_din )
       end
endmodule // gdp

`ifdef TEST
module test ;

   parameter W = 32 ;//Width of data input bus
   parameter N = 3 ;//Number of data words in packet
   parameter LOG2N = 2 ;//Ceiling of Log2(N)
   
   parameter BIGENDIAN = 0;//1 if big endian

   /*AUTOREGINPUT*/
   // Beginning of automatic reg inputs (for undeclared instantiated-module inputs)
   reg			clk;			// To dut of gdu.v
   reg [W-1:0]		din;			// To dut of gdu.v
   reg			eop;			// To dut of gdu.v
   reg			reset;			// To dut of gdu.v
   reg			sop;			// To dut of gdu.v
   reg			valid_din;		// To dut of gdu.v
   // End of automatics

   /*AUTOWIRE*/
   // Beginning of automatic wires (for undeclared instantiated-module outputs)
   wire [`F0_W-1:0]	dout_f0;		// From dut of gdu.v
   wire [`F1_W-1:0]	dout_f1;		// From dut of gdu.v
   wire [`F2_W-1:0]	dout_f2;		// From dut of gdu.v
   wire [`F3_W-1:0]	dout_f3;		// From dut of gdu.v
   wire [`F4_W-1:0]	dout_f4;		// From dut of gdu.v
   wire			err;			// From dut of gdu.v
   wire			valid_f0;		// From dut of gdu.v
   wire			valid_f1;		// From dut of gdu.v
   wire			valid_f2;		// From dut of gdu.v
   wire			valid_f3;		// From dut of gdu.v
   wire			valid_f4;		// From dut of gdu.v
   // End of automatics
   
   initial
     begin
	$dumpvars;
	clk = 0;
	din = 0;
	eop = 0;
	sop = 0;
	reset = 0;
	valid_din = 0;
	reset_dut;
	repeat(20) $display("random no = %d",$random);
       	repeat (20000) @(posedge clk);
	$finish;
     end

   always #5 clk = ~clk ;

   task reset_dut;
     begin
	@(posedge clk);
	reset <= 1;
	repeat (20) @(posedge clk);
	reset <= 0;
	repeat (20) @(posedge clk);	
     end
   endtask // reset_dut

   always @(posedge clk)
     begin
	if ($random % 4)
	  begin
	     din <= din + 1;
	     valid_din <= 1;
	  end
	else
	  valid_din <= 0;
     end

   gdu dut (/*AUTOINST*/
	    // Outputs
	    .err			(err),
	    .valid_f0			(valid_f0),
	    .valid_f1			(valid_f1),
	    .valid_f2			(valid_f2),
	    .valid_f3			(valid_f3),
	    .valid_f4			(valid_f4),
	    .dout_f0			(dout_f0[`F0_W-1:0]),
	    .dout_f1			(dout_f1[`F1_W-1:0]),
	    .dout_f2			(dout_f2[`F2_W-1:0]),
	    .dout_f3			(dout_f3[`F3_W-1:0]),
	    .dout_f4			(dout_f4[`F4_W-1:0]),
	    // Inputs
	    .clk			(clk),
	    .reset			(reset),
	    .sop			(sop),
	    .eop			(eop),
	    .din			(din[W-1:0]),
	    .valid_din			(valid_din));
   

endmodule  // test

`endif

