`define f0_W0_LSB  0
`define f0_W0_MSB  4

`define f1_W0_LSB  5
`define f1_W0_MSB  10

`define f2_W0_LSB  11
`define f2_W0_MSB  31
`define f2_W1_LSB  0
`define f2_W1_MSB  40

`define f3_W1_LSB  41
`define f3_W1_MSB  31
`define f3_W2_LSB  0
`define f3_W2_MSB  13

`define f4_W2_LSB  14
`define f4_W2_MSB  31
`define f4_W3_LSB  0
`define f4_W3_MSB  4

`define f5_W3_LSB  5
`define f5_W3_MSB  31
`define f5_W4_LSB  0
`define f5_W4_MSB  4

`define f6_W4_LSB  5
`define f6_W4_MSB  27

`define f7_W4_LSB  28
`define f7_W4_MSB  31
`define f7_W5_LSB  0
`define f7_W5_MSB  1

`define f8_W5_LSB  2
`define f8_W5_MSB  31
`define f8_W6_LSB  0
`define f8_W6_MSB  1

`define f9_W6_LSB  2
`define f9_W6_MSB  31

