`timescale 1ns/1ps

`define ENABLED_REGEX_ALL_0 TRUE

module ALL_0_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_ALL_0

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd8;
    1: charMap = 8'd8;
    2: charMap = 8'd8;
    3: charMap = 8'd8;
    4: charMap = 8'd8;
    5: charMap = 8'd8;
    6: charMap = 8'd8;
    7: charMap = 8'd8;
    8: charMap = 8'd8;
    9: charMap = 8'd20;
    10: charMap = 8'd21;
    11: charMap = 8'd20;
    12: charMap = 8'd8;
    13: charMap = 8'd21;
    14: charMap = 8'd8;
    15: charMap = 8'd8;
    16: charMap = 8'd8;
    17: charMap = 8'd8;
    18: charMap = 8'd8;
    19: charMap = 8'd8;
    20: charMap = 8'd8;
    21: charMap = 8'd8;
    22: charMap = 8'd8;
    23: charMap = 8'd8;
    24: charMap = 8'd8;
    25: charMap = 8'd8;
    26: charMap = 8'd8;
    27: charMap = 8'd8;
    28: charMap = 8'd8;
    29: charMap = 8'd8;
    30: charMap = 8'd8;
    31: charMap = 8'd8;
    32: charMap = 8'd20;
    33: charMap = 8'd8;
    34: charMap = 8'd23;
    35: charMap = 8'd8;
    36: charMap = 8'd8;
    37: charMap = 8'd29;
    38: charMap = 8'd25;
    39: charMap = 8'd24;
    40: charMap = 8'd22;
    41: charMap = 8'd8;
    42: charMap = 8'd8;
    43: charMap = 8'd31;
    44: charMap = 8'd8;
    45: charMap = 8'd8;
    46: charMap = 8'd8;
    47: charMap = 8'd8;
    48: charMap = 8'd30;
    49: charMap = 8'd30;
    50: charMap = 8'd30;
    51: charMap = 8'd30;
    52: charMap = 8'd30;
    53: charMap = 8'd30;
    54: charMap = 8'd30;
    55: charMap = 8'd30;
    56: charMap = 8'd30;
    57: charMap = 8'd30;
    58: charMap = 8'd8;
    59: charMap = 8'd27;
    60: charMap = 8'd8;
    61: charMap = 8'd8;
    62: charMap = 8'd8;
    63: charMap = 8'd8;
    64: charMap = 8'd8;
    65: charMap = 8'd8;
    66: charMap = 8'd8;
    67: charMap = 8'd8;
    68: charMap = 8'd8;
    69: charMap = 8'd8;
    70: charMap = 8'd8;
    71: charMap = 8'd8;
    72: charMap = 8'd8;
    73: charMap = 8'd8;
    74: charMap = 8'd8;
    75: charMap = 8'd8;
    76: charMap = 8'd8;
    77: charMap = 8'd8;
    78: charMap = 8'd8;
    79: charMap = 8'd8;
    80: charMap = 8'd8;
    81: charMap = 8'd8;
    82: charMap = 8'd8;
    83: charMap = 8'd8;
    84: charMap = 8'd8;
    85: charMap = 8'd8;
    86: charMap = 8'd8;
    87: charMap = 8'd8;
    88: charMap = 8'd8;
    89: charMap = 8'd8;
    90: charMap = 8'd8;
    91: charMap = 8'd8;
    92: charMap = 8'd28;
    93: charMap = 8'd8;
    94: charMap = 8'd8;
    95: charMap = 8'd12;
    96: charMap = 8'd8;
    97: charMap = 8'd6;
    98: charMap = 8'd17;
    99: charMap = 8'd5;
    100: charMap = 8'd13;
    101: charMap = 8'd3;
    102: charMap = 8'd30;
    103: charMap = 8'd19;
    104: charMap = 8'd16;
    105: charMap = 8'd8;
    106: charMap = 8'd8;
    107: charMap = 8'd18;
    108: charMap = 8'd14;
    109: charMap = 8'd8;
    110: charMap = 8'd2;
    111: charMap = 8'd15;
    112: charMap = 8'd7;
    113: charMap = 8'd26;
    114: charMap = 8'd9;
    115: charMap = 8'd4;
    116: charMap = 8'd11;
    117: charMap = 8'd1;
    118: charMap = 8'd8;
    119: charMap = 8'd8;
    120: charMap = 8'd8;
    121: charMap = 8'd10;
    122: charMap = 8'd8;
    123: charMap = 8'd8;
    124: charMap = 8'd8;
    125: charMap = 8'd8;
    126: charMap = 8'd8;
    127: charMap = 8'd8;
    128: charMap = 8'd8;
    129: charMap = 8'd8;
    130: charMap = 8'd8;
    131: charMap = 8'd8;
    132: charMap = 8'd8;
    133: charMap = 8'd8;
    134: charMap = 8'd8;
    135: charMap = 8'd8;
    136: charMap = 8'd8;
    137: charMap = 8'd8;
    138: charMap = 8'd8;
    139: charMap = 8'd8;
    140: charMap = 8'd8;
    141: charMap = 8'd8;
    142: charMap = 8'd8;
    143: charMap = 8'd8;
    144: charMap = 8'd8;
    145: charMap = 8'd8;
    146: charMap = 8'd8;
    147: charMap = 8'd8;
    148: charMap = 8'd8;
    149: charMap = 8'd8;
    150: charMap = 8'd8;
    151: charMap = 8'd8;
    152: charMap = 8'd8;
    153: charMap = 8'd8;
    154: charMap = 8'd8;
    155: charMap = 8'd8;
    156: charMap = 8'd8;
    157: charMap = 8'd8;
    158: charMap = 8'd8;
    159: charMap = 8'd8;
    160: charMap = 8'd8;
    161: charMap = 8'd8;
    162: charMap = 8'd8;
    163: charMap = 8'd8;
    164: charMap = 8'd8;
    165: charMap = 8'd8;
    166: charMap = 8'd8;
    167: charMap = 8'd8;
    168: charMap = 8'd8;
    169: charMap = 8'd8;
    170: charMap = 8'd8;
    171: charMap = 8'd8;
    172: charMap = 8'd8;
    173: charMap = 8'd8;
    174: charMap = 8'd8;
    175: charMap = 8'd8;
    176: charMap = 8'd8;
    177: charMap = 8'd8;
    178: charMap = 8'd8;
    179: charMap = 8'd8;
    180: charMap = 8'd8;
    181: charMap = 8'd8;
    182: charMap = 8'd8;
    183: charMap = 8'd8;
    184: charMap = 8'd8;
    185: charMap = 8'd8;
    186: charMap = 8'd8;
    187: charMap = 8'd8;
    188: charMap = 8'd8;
    189: charMap = 8'd8;
    190: charMap = 8'd8;
    191: charMap = 8'd8;
    192: charMap = 8'd8;
    193: charMap = 8'd8;
    194: charMap = 8'd8;
    195: charMap = 8'd8;
    196: charMap = 8'd8;
    197: charMap = 8'd8;
    198: charMap = 8'd8;
    199: charMap = 8'd8;
    200: charMap = 8'd8;
    201: charMap = 8'd8;
    202: charMap = 8'd8;
    203: charMap = 8'd8;
    204: charMap = 8'd8;
    205: charMap = 8'd8;
    206: charMap = 8'd8;
    207: charMap = 8'd8;
    208: charMap = 8'd8;
    209: charMap = 8'd8;
    210: charMap = 8'd8;
    211: charMap = 8'd8;
    212: charMap = 8'd8;
    213: charMap = 8'd8;
    214: charMap = 8'd8;
    215: charMap = 8'd8;
    216: charMap = 8'd8;
    217: charMap = 8'd8;
    218: charMap = 8'd8;
    219: charMap = 8'd8;
    220: charMap = 8'd8;
    221: charMap = 8'd8;
    222: charMap = 8'd8;
    223: charMap = 8'd8;
    224: charMap = 8'd8;
    225: charMap = 8'd8;
    226: charMap = 8'd8;
    227: charMap = 8'd8;
    228: charMap = 8'd8;
    229: charMap = 8'd8;
    230: charMap = 8'd8;
    231: charMap = 8'd8;
    232: charMap = 8'd8;
    233: charMap = 8'd8;
    234: charMap = 8'd8;
    235: charMap = 8'd8;
    236: charMap = 8'd8;
    237: charMap = 8'd8;
    238: charMap = 8'd8;
    239: charMap = 8'd8;
    240: charMap = 8'd8;
    241: charMap = 8'd8;
    242: charMap = 8'd8;
    243: charMap = 8'd8;
    244: charMap = 8'd8;
    245: charMap = 8'd8;
    246: charMap = 8'd8;
    247: charMap = 8'd8;
    248: charMap = 8'd8;
    249: charMap = 8'd8;
    250: charMap = 8'd8;
    251: charMap = 8'd8;
    252: charMap = 8'd8;
    253: charMap = 8'd8;
    254: charMap = 8'd8;
    255: charMap = 8'd8;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd2;
    3: stateMap = 11'd3;
    4: stateMap = 11'd1;
    5: stateMap = 11'd4;
    6: stateMap = 11'd5;
    7: stateMap = 11'd6;
    8: stateMap = 11'd7;
    9: stateMap = 11'd8;
    10: stateMap = 11'd9;
    11: stateMap = 11'd10;
    12: stateMap = 11'd11;
    13: stateMap = 11'd12;
    14: stateMap = 11'd13;
    15: stateMap = 11'd14;
    16: stateMap = 11'd15;
    17: stateMap = 11'd16;
    18: stateMap = 11'd17;
    19: stateMap = 11'd18;
    20: stateMap = 11'd19;
    21: stateMap = 11'd20;
    22: stateMap = 11'd21;
    23: stateMap = 11'd22;
    24: stateMap = 11'd23;
    25: stateMap = 11'd24;
    26: stateMap = 11'd25;
    27: stateMap = 11'd26;
    28: stateMap = 11'd27;
    29: stateMap = 11'd28;
    30: stateMap = 11'd29;
    31: stateMap = 11'd30;
    32: stateMap = 11'd31;
    33: stateMap = 11'd32;
    34: stateMap = 11'd33;
    35: stateMap = 11'd34;
    36: stateMap = 11'd35;
    37: stateMap = 11'd36;
    38: stateMap = 11'd37;
    39: stateMap = 11'd38;
    40: stateMap = 11'd39;
    41: stateMap = 11'd40;
    42: stateMap = 11'd41;
    43: stateMap = 11'd42;
    44: stateMap = 11'd43;
    45: stateMap = 11'd44;
    46: stateMap = 11'd45;
    47: stateMap = 11'd46;
    48: stateMap = 11'd47;
    49: stateMap = 11'd48;
    50: stateMap = 11'd49;
    51: stateMap = 11'd50;
    52: stateMap = 11'd51;
    53: stateMap = 11'd52;
    54: stateMap = 11'd53;
    55: stateMap = 11'd54;
    56: stateMap = 11'd55;
    57: stateMap = 11'd56;
    58: stateMap = 11'd57;
    59: stateMap = 11'd2;
    60: stateMap = 11'd58;
    61: stateMap = 11'd59;
    62: stateMap = 11'd60;
    63: stateMap = 11'd56;
    64: stateMap = 11'd61;
    65: stateMap = 11'd62;
    66: stateMap = 11'd2;
    67: stateMap = 11'd63;
    68: stateMap = 11'd64;
    69: stateMap = 11'd60;
    70: stateMap = 11'd65;
    71: stateMap = 11'd66;
    72: stateMap = 11'd67;
    73: stateMap = 11'd68;
    74: stateMap = 11'd69;
    75: stateMap = 11'd70;
    76: stateMap = 11'd71;
    77: stateMap = 11'd72;
    78: stateMap = 11'd73;
    79: stateMap = 11'd74;
    80: stateMap = 11'd75;
    81: stateMap = 11'd76;
    82: stateMap = 11'd66;
    83: stateMap = 11'd77;
    84: stateMap = 11'd78;
    85: stateMap = 11'd68;
    86: stateMap = 11'd79;
    87: stateMap = 11'd80;
    88: stateMap = 11'd81;
    89: stateMap = 11'd82;
    90: stateMap = 11'd83;
    91: stateMap = 11'd84;
    92: stateMap = 11'd85;
    93: stateMap = 11'd86;
    94: stateMap = 11'd87;
    95: stateMap = 11'd88;
    96: stateMap = 11'd82;
    97: stateMap = 11'd89;
    98: stateMap = 11'd86;
    99: stateMap = 11'd90;
    100: stateMap = 11'd91;
    101: stateMap = 11'd92;
    102: stateMap = 11'd93;
    103: stateMap = 11'd94;
    104: stateMap = 11'd95;
    105: stateMap = 11'd96;
    106: stateMap = 11'd97;
    107: stateMap = 11'd98;
    108: stateMap = 11'd99;
    109: stateMap = 11'd100;
    110: stateMap = 11'd101;
    111: stateMap = 11'd102;
    112: stateMap = 11'd103;
    113: stateMap = 11'd104;
    114: stateMap = 11'd105;
    115: stateMap = 11'd106;
    116: stateMap = 11'd107;
    117: stateMap = 11'd108;
    118: stateMap = 11'd109;
    119: stateMap = 11'd110;
    120: stateMap = 11'd111;
    121: stateMap = 11'd112;
    122: stateMap = 11'd113;
    123: stateMap = 11'd114;
    124: stateMap = 11'd115;
    125: stateMap = 11'd116;
    126: stateMap = 11'd117;
    127: stateMap = 11'd118;
    128: stateMap = 11'd119;
    129: stateMap = 11'd120;
    130: stateMap = 11'd121;
    131: stateMap = 11'd122;
    132: stateMap = 11'd123;
    133: stateMap = 11'd124;
    134: stateMap = 11'd125;
    135: stateMap = 11'd126;
    136: stateMap = 11'd127;
    137: stateMap = 11'd128;
    138: stateMap = 11'd129;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b1;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b0;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b0;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b0;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b0;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b0;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b0;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b0;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b0;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b0;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b0;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b0;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b0;
    62: acceptStates = 1'b0;
    63: acceptStates = 1'b0;
    64: acceptStates = 1'b0;
    65: acceptStates = 1'b0;
    66: acceptStates = 1'b0;
    67: acceptStates = 1'b0;
    68: acceptStates = 1'b0;
    69: acceptStates = 1'b0;
    70: acceptStates = 1'b0;
    71: acceptStates = 1'b0;
    72: acceptStates = 1'b0;
    73: acceptStates = 1'b0;
    74: acceptStates = 1'b0;
    75: acceptStates = 1'b0;
    76: acceptStates = 1'b0;
    77: acceptStates = 1'b0;
    78: acceptStates = 1'b0;
    79: acceptStates = 1'b0;
    80: acceptStates = 1'b0;
    81: acceptStates = 1'b0;
    82: acceptStates = 1'b0;
    83: acceptStates = 1'b0;
    84: acceptStates = 1'b0;
    85: acceptStates = 1'b0;
    86: acceptStates = 1'b0;
    87: acceptStates = 1'b0;
    88: acceptStates = 1'b0;
    89: acceptStates = 1'b0;
    90: acceptStates = 1'b0;
    91: acceptStates = 1'b0;
    92: acceptStates = 1'b0;
    93: acceptStates = 1'b0;
    94: acceptStates = 1'b0;
    95: acceptStates = 1'b0;
    96: acceptStates = 1'b0;
    97: acceptStates = 1'b0;
    98: acceptStates = 1'b0;
    99: acceptStates = 1'b0;
    100: acceptStates = 1'b0;
    101: acceptStates = 1'b0;
    102: acceptStates = 1'b0;
    103: acceptStates = 1'b0;
    104: acceptStates = 1'b0;
    105: acceptStates = 1'b0;
    106: acceptStates = 1'b0;
    107: acceptStates = 1'b0;
    108: acceptStates = 1'b0;
    109: acceptStates = 1'b0;
    110: acceptStates = 1'b0;
    111: acceptStates = 1'b0;
    112: acceptStates = 1'b0;
    113: acceptStates = 1'b0;
    114: acceptStates = 1'b0;
    115: acceptStates = 1'b0;
    116: acceptStates = 1'b0;
    117: acceptStates = 1'b0;
    118: acceptStates = 1'b0;
    119: acceptStates = 1'b0;
    120: acceptStates = 1'b0;
    121: acceptStates = 1'b0;
    122: acceptStates = 1'b0;
    123: acceptStates = 1'b0;
    124: acceptStates = 1'b0;
    125: acceptStates = 1'b0;
    126: acceptStates = 1'b0;
    127: acceptStates = 1'b0;
    128: acceptStates = 1'b0;
    129: acceptStates = 1'b0;
    130: acceptStates = 1'b0;
    131: acceptStates = 1'b0;
    132: acceptStates = 1'b0;
    133: acceptStates = 1'b0;
    134: acceptStates = 1'b0;
    135: acceptStates = 1'b0;
    136: acceptStates = 1'b0;
    137: acceptStates = 1'b0;
    138: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd1;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd5;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd6;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd7;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd8;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd9;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd10;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd12;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd77;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd13;
      21: stateTransition = 11'd13;
      22: stateTransition = 11'd14;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd15;
      24: stateTransition = 11'd15;
      25: stateTransition = 11'd16;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd17;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd18;
      29: stateTransition = 11'd18;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd33;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd15;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd44;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd44;
      6: stateTransition = 11'd44;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd44;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd44;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd44;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd21;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd22;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd15;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd25;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd26;
      29: stateTransition = 11'd26;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd24;
      21: stateTransition = 11'd25;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd27;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd25;
      21: stateTransition = 11'd25;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd28;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd46;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd27;
      21: stateTransition = 11'd28;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd51;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd28;
      21: stateTransition = 11'd28;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd32;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd2;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd2;
      6: stateTransition = 11'd2;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd2;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd2;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd2;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd4;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd4;
      6: stateTransition = 11'd4;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd4;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd4;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd4;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd12;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd26;
      29: stateTransition = 11'd26;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd20;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd0;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd23;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd23;
      6: stateTransition = 11'd23;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd23;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd23;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd23;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd24;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd50;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd30;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd30;
      6: stateTransition = 11'd30;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd30;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd30;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd30;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd29;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd29;
      6: stateTransition = 11'd29;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd29;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd29;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd29;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd31;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd34;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd34;
      6: stateTransition = 11'd34;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd34;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd34;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd34;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd35;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd35;
      6: stateTransition = 11'd35;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd35;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd35;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd35;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd36;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd36;
      6: stateTransition = 11'd36;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd36;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd36;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd36;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd37;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd37;
      6: stateTransition = 11'd37;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd37;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd37;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd37;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd38;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd39;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd39;
      6: stateTransition = 11'd39;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd39;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd39;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd39;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd40;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd40;
      6: stateTransition = 11'd40;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd40;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd40;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd40;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd41;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd41;
      6: stateTransition = 11'd41;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd41;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd41;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      30: stateTransition = 11'd41;
      31: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd42;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd42;
      6: stateTransition = 11'd42;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd42;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd42;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd42;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd43;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd85;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd45;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd45;
      6: stateTransition = 11'd45;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd45;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd45;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd45;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd47;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd50;
      29: stateTransition = 11'd50;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd48;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd49;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd49;
      6: stateTransition = 11'd49;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd49;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd49;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd49;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd52;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd134;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd53;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd56;
      29: stateTransition = 11'd56;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd55;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd105;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd89;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd60;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    60: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd61;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    61: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd57;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    62: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd57;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    63: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd60;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    64: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    65: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd116;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    66: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd67;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    67: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd69;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    68: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd71;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    69: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    70: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd62;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    71: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd93;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd115;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd135;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    72: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd63;
      24: stateTransition = 11'd63;
      25: stateTransition = 11'd78;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd64;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    73: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd83;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    74: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd65;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    75: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd117;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd104;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd66;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    76: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd79;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    77: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd81;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    78: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd68;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    79: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd66;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd116;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    80: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd73;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    81: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd70;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    82: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd93;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd85;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    83: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd72;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    84: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd75;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    85: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd74;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    86: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd85;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    87: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd76;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd119;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    88: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd100;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    89: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd80;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd135;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    90: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd96;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd60;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    91: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd99;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    92: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd66;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    93: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd84;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    94: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd87;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    95: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd127;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd86;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    96: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd91;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    97: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd101;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    98: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd95;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    99: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd88;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    100: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd90;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd116;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    101: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd92;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    102: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd94;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    103: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd97;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    104: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd107;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    105: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd102;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    106: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd117;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd104;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    107: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd106;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    108: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd118;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd116;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    109: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd108;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    110: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd137;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd109;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    111: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd110;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    112: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd131;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd116;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    113: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd111;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    114: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd115;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd135;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    115: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd113;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    116: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd116;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    117: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd117;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    118: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd119;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    119: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd120;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    120: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd138;
      3: stateTransition = 11'd127;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    121: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd121;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    122: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd122;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    123: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd127;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    124: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd59;
      3: stateTransition = 11'd59;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd124;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    125: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd58;
      2: stateTransition = 11'd133;
      3: stateTransition = 11'd67;
      4: stateTransition = 11'd98;
      5: stateTransition = 11'd59;
      6: stateTransition = 11'd59;
      7: stateTransition = 11'd59;
      8: stateTransition = 11'd59;
      9: stateTransition = 11'd82;
      10: stateTransition = 11'd59;
      11: stateTransition = 11'd59;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd59;
      14: stateTransition = 11'd59;
      15: stateTransition = 11'd59;
      16: stateTransition = 11'd103;
      17: stateTransition = 11'd59;
      18: stateTransition = 11'd59;
      19: stateTransition = 11'd59;
      20: stateTransition = 11'd59;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd59;
      23: stateTransition = 11'd59;
      24: stateTransition = 11'd59;
      25: stateTransition = 11'd59;
      26: stateTransition = 11'd59;
      27: stateTransition = 11'd59;
      28: stateTransition = 11'd59;
      29: stateTransition = 11'd59;
      30: stateTransition = 11'd59;
      31: stateTransition = 11'd59;
      default: stateTransition = 11'bX;
    endcase
    126: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd136;
      4: stateTransition = 11'd97;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    127: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd128;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    128: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd129;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd11;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    129: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd11;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd11;
      4: stateTransition = 11'd123;
      5: stateTransition = 11'd11;
      6: stateTransition = 11'd125;
      7: stateTransition = 11'd126;
      8: stateTransition = 11'd11;
      9: stateTransition = 11'd132;
      10: stateTransition = 11'd11;
      11: stateTransition = 11'd11;
      12: stateTransition = 11'd130;
      13: stateTransition = 11'd11;
      14: stateTransition = 11'd11;
      15: stateTransition = 11'd11;
      16: stateTransition = 11'd112;
      17: stateTransition = 11'd114;
      18: stateTransition = 11'd11;
      19: stateTransition = 11'd11;
      20: stateTransition = 11'd11;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd11;
      23: stateTransition = 11'd11;
      24: stateTransition = 11'd11;
      25: stateTransition = 11'd11;
      26: stateTransition = 11'd11;
      27: stateTransition = 11'd11;
      28: stateTransition = 11'd11;
      29: stateTransition = 11'd11;
      30: stateTransition = 11'd11;
      31: stateTransition = 11'd11;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
