wire fired_ALL_0 ;
wire fired_ALL_10 ;
wire fired_ALL_11 ;
wire fired_ALL_12 ;
wire fired_ALL_13 ;
wire fired_ALL_14 ;
wire fired_ALL_1 ;
wire fired_ALL_2 ;
wire fired_ALL_3 ;
wire fired_ALL_4 ;
wire fired_ALL_5 ;
wire fired_ALL_6 ;
wire fired_ALL_7 ;
wire fired_ALL_8 ;
wire fired_ALL_9 ;
wire fired_finger_0 ;
wire fired_finger_1 ;
wire fired_finger_2 ;
wire fired_finger_3 ;
wire fired_finger_4 ;
wire fired_finger_5 ;
wire fired_ftp_0 ;
wire fired_ftp_1 ;
wire fired_ftp_2 ;
wire fired_ftp_3 ;
wire fired_ftp_4 ;
wire fired_ftp_5 ;
wire fired_ftp_6 ;
wire fired_ftp_7 ;
wire fired_ftp_8 ;
wire fired_ftp_9 ;
wire fired_http_0 ;
wire fired_http_1 ;
wire fired_http_2 ;
wire fired_http_3 ;
wire fired_http_4 ;
wire fired_http_5 ;
wire fired_http_6 ;
wire fired_http_7 ;
wire fired_http_8 ;
wire fired_http_9 ;
wire fired_imap_0 ;
wire fired_imap_1 ;
wire fired_imap_2 ;
wire fired_imap_3 ;
wire fired_imap_4 ;
wire fired_imap_5 ;
wire fired_imap_6 ;
wire fired_imap_7 ;
wire fired_imap_8 ;
wire fired_imap_9 ;
wire fired_netbios_0 ;
wire fired_netbios_1 ;
wire fired_netbios_2 ;
wire fired_netbios_3 ;
wire fired_netbios_4 ;
wire fired_netbios_5 ;
wire fired_netbios_6 ;
wire fired_netbios_7 ;
wire fired_netbios_8 ;
wire fired_netbios_9 ;
wire fired_nntp_0 ;
wire fired_nntp_1 ;
wire fired_nntp_2 ;
wire fired_nntp_3 ;
wire fired_nntp_4 ;
wire fired_nntp_5 ;
wire fired_nntp_6 ;
wire fired_nntp_7 ;
wire fired_nntp_8 ;
wire fired_nntp_9 ;
wire fired_pop3_0 ;
wire fired_pop3_1 ;
wire fired_pop3_2 ;
wire fired_pop3_3 ;
wire fired_pop3_4 ;
wire fired_pop3_5 ;
wire fired_pop3_6 ;
wire fired_pop3_7 ;
wire fired_pop3_8 ;
wire fired_pop3_9 ;
wire fired_rlogin_0 ;
wire fired_rlogin_1 ;
wire fired_rlogin_2 ;
wire fired_rlogin_3 ;
wire fired_rlogin_4 ;
wire fired_rlogin_5 ;
wire fired_smtp_0 ;
wire fired_smtp_1 ;
wire fired_smtp_2 ;
wire fired_smtp_3 ;
wire fired_smtp_4 ;
wire fired_smtp_5 ;
wire fired_smtp_6 ;
wire fired_smtp_7 ;
wire fired_smtp_8 ;
wire fired_smtp_9 ;
wire fired_telnet_0 ;
wire fired_telnet_1 ;
wire fired_telnet_2 ;
wire fired_telnet_3 ;
wire fired_telnet_4 ;
wire fired_telnet_5 ;
wire fired_telnet_6 ;
wire fired_telnet_7 ;
wire fired_telnet_8 ;
wire fired_telnet_9 ;
wire fired_CATEGORY_aim ;
wire fired_CATEGORY_bittorrent ;
wire fired_CATEGORY_cvs ;
wire fired_CATEGORY_dhcp ;
wire fired_CATEGORY_directconnect ;
wire fired_CATEGORY_dns ;
wire fired_CATEGORY_fasttrack ;
wire fired_CATEGORY_finger ;
wire fired_CATEGORY_freenet ;
wire fired_CATEGORY_ftp ;
wire fired_CATEGORY_gnutella ;
wire fired_CATEGORY_gopher ;
wire fired_CATEGORY_http ;
wire fired_CATEGORY_imap ;
wire fired_CATEGORY_irc ;
wire fired_CATEGORY_jabber ;
wire fired_CATEGORY_msn ;
wire fired_CATEGORY_napster ;
wire fired_CATEGORY_netbios ;
wire fired_CATEGORY_nntp ;
wire fired_CATEGORY_pop3 ;
wire fired_CATEGORY_rlogin ;
wire fired_CATEGORY_sip ;
wire fired_CATEGORY_smtp ;
wire fired_CATEGORY_snmp ;
wire fired_CATEGORY_socks ;
wire fired_CATEGORY_ssh ;
wire fired_CATEGORY_ssl ;
wire fired_CATEGORY_subversion ;
wire fired_CATEGORY_telnet ;
wire fired_CATEGORY_tor ;
wire fired_CATEGORY_vnc ;
wire fired_CATEGORY_worldofwarcraft ;
wire fired_CATEGORY_x11 ;
wire fired_CATEGORY_yahoo ;
