`timescale 1ns/1ps

`define ENABLED_REGEX_ALL_3 TRUE

module ALL_3_verilog(clk,
                    rst_n,
                    char_in,
                    char_in_vld,
                    state_in,
                    state_in_vld,
                    state_out,
                    accept_out);
   // The clock and reset info.
    input clk, rst_n;
    // Input character, and state, if being set.
    input [7:0] char_in;
    input [10:0] state_in;
    // char_in_vld should be true if there's a character to process.
    // state_in_vld should be true if the outside world is overwriting our state.
    input char_in_vld, state_in_vld;
    // state_out is our current state.
    output [10:0] state_out;
    // Accept out is true if the character triggered a regex match.
    output accept_out;
    // A register for the current state.
    reg [10:0] cur_state;


`ifdef ENABLED_REGEX_ALL_3

function [7:0] charMap;
  input [7:0] inchar;
  begin
  case( inchar )
    0: charMap = 8'd2;
    1: charMap = 8'd9;
    2: charMap = 8'd9;
    3: charMap = 8'd9;
    4: charMap = 8'd9;
    5: charMap = 8'd9;
    6: charMap = 8'd9;
    7: charMap = 8'd9;
    8: charMap = 8'd9;
    9: charMap = 8'd21;
    10: charMap = 8'd22;
    11: charMap = 8'd21;
    12: charMap = 8'd9;
    13: charMap = 8'd22;
    14: charMap = 8'd9;
    15: charMap = 8'd9;
    16: charMap = 8'd9;
    17: charMap = 8'd9;
    18: charMap = 8'd9;
    19: charMap = 8'd9;
    20: charMap = 8'd9;
    21: charMap = 8'd9;
    22: charMap = 8'd9;
    23: charMap = 8'd9;
    24: charMap = 8'd9;
    25: charMap = 8'd9;
    26: charMap = 8'd9;
    27: charMap = 8'd9;
    28: charMap = 8'd9;
    29: charMap = 8'd9;
    30: charMap = 8'd9;
    31: charMap = 8'd9;
    32: charMap = 8'd21;
    33: charMap = 8'd9;
    34: charMap = 8'd24;
    35: charMap = 8'd9;
    36: charMap = 8'd9;
    37: charMap = 8'd9;
    38: charMap = 8'd26;
    39: charMap = 8'd25;
    40: charMap = 8'd23;
    41: charMap = 8'd9;
    42: charMap = 8'd9;
    43: charMap = 8'd9;
    44: charMap = 8'd9;
    45: charMap = 8'd9;
    46: charMap = 8'd9;
    47: charMap = 8'd9;
    48: charMap = 8'd9;
    49: charMap = 8'd9;
    50: charMap = 8'd9;
    51: charMap = 8'd9;
    52: charMap = 8'd9;
    53: charMap = 8'd9;
    54: charMap = 8'd9;
    55: charMap = 8'd9;
    56: charMap = 8'd9;
    57: charMap = 8'd9;
    58: charMap = 8'd9;
    59: charMap = 8'd28;
    60: charMap = 8'd9;
    61: charMap = 8'd9;
    62: charMap = 8'd9;
    63: charMap = 8'd9;
    64: charMap = 8'd9;
    65: charMap = 8'd9;
    66: charMap = 8'd9;
    67: charMap = 8'd9;
    68: charMap = 8'd9;
    69: charMap = 8'd9;
    70: charMap = 8'd9;
    71: charMap = 8'd9;
    72: charMap = 8'd9;
    73: charMap = 8'd9;
    74: charMap = 8'd9;
    75: charMap = 8'd9;
    76: charMap = 8'd9;
    77: charMap = 8'd9;
    78: charMap = 8'd9;
    79: charMap = 8'd9;
    80: charMap = 8'd9;
    81: charMap = 8'd9;
    82: charMap = 8'd9;
    83: charMap = 8'd9;
    84: charMap = 8'd9;
    85: charMap = 8'd9;
    86: charMap = 8'd9;
    87: charMap = 8'd9;
    88: charMap = 8'd9;
    89: charMap = 8'd9;
    90: charMap = 8'd9;
    91: charMap = 8'd9;
    92: charMap = 8'd29;
    93: charMap = 8'd9;
    94: charMap = 8'd9;
    95: charMap = 8'd13;
    96: charMap = 8'd9;
    97: charMap = 8'd7;
    98: charMap = 8'd18;
    99: charMap = 8'd6;
    100: charMap = 8'd14;
    101: charMap = 8'd4;
    102: charMap = 8'd9;
    103: charMap = 8'd20;
    104: charMap = 8'd17;
    105: charMap = 8'd9;
    106: charMap = 8'd9;
    107: charMap = 8'd19;
    108: charMap = 8'd15;
    109: charMap = 8'd9;
    110: charMap = 8'd3;
    111: charMap = 8'd16;
    112: charMap = 8'd8;
    113: charMap = 8'd27;
    114: charMap = 8'd10;
    115: charMap = 8'd5;
    116: charMap = 8'd12;
    117: charMap = 8'd1;
    118: charMap = 8'd9;
    119: charMap = 8'd9;
    120: charMap = 8'd9;
    121: charMap = 8'd11;
    122: charMap = 8'd9;
    123: charMap = 8'd9;
    124: charMap = 8'd9;
    125: charMap = 8'd9;
    126: charMap = 8'd9;
    127: charMap = 8'd9;
    128: charMap = 8'd9;
    129: charMap = 8'd9;
    130: charMap = 8'd9;
    131: charMap = 8'd9;
    132: charMap = 8'd9;
    133: charMap = 8'd9;
    134: charMap = 8'd9;
    135: charMap = 8'd9;
    136: charMap = 8'd9;
    137: charMap = 8'd9;
    138: charMap = 8'd9;
    139: charMap = 8'd9;
    140: charMap = 8'd9;
    141: charMap = 8'd9;
    142: charMap = 8'd9;
    143: charMap = 8'd9;
    144: charMap = 8'd9;
    145: charMap = 8'd9;
    146: charMap = 8'd9;
    147: charMap = 8'd9;
    148: charMap = 8'd9;
    149: charMap = 8'd9;
    150: charMap = 8'd9;
    151: charMap = 8'd9;
    152: charMap = 8'd9;
    153: charMap = 8'd9;
    154: charMap = 8'd9;
    155: charMap = 8'd9;
    156: charMap = 8'd9;
    157: charMap = 8'd9;
    158: charMap = 8'd9;
    159: charMap = 8'd9;
    160: charMap = 8'd9;
    161: charMap = 8'd9;
    162: charMap = 8'd9;
    163: charMap = 8'd9;
    164: charMap = 8'd9;
    165: charMap = 8'd9;
    166: charMap = 8'd9;
    167: charMap = 8'd9;
    168: charMap = 8'd9;
    169: charMap = 8'd9;
    170: charMap = 8'd9;
    171: charMap = 8'd9;
    172: charMap = 8'd9;
    173: charMap = 8'd9;
    174: charMap = 8'd9;
    175: charMap = 8'd9;
    176: charMap = 8'd9;
    177: charMap = 8'd9;
    178: charMap = 8'd9;
    179: charMap = 8'd9;
    180: charMap = 8'd9;
    181: charMap = 8'd9;
    182: charMap = 8'd9;
    183: charMap = 8'd9;
    184: charMap = 8'd9;
    185: charMap = 8'd9;
    186: charMap = 8'd9;
    187: charMap = 8'd9;
    188: charMap = 8'd9;
    189: charMap = 8'd9;
    190: charMap = 8'd9;
    191: charMap = 8'd9;
    192: charMap = 8'd9;
    193: charMap = 8'd9;
    194: charMap = 8'd9;
    195: charMap = 8'd9;
    196: charMap = 8'd9;
    197: charMap = 8'd9;
    198: charMap = 8'd9;
    199: charMap = 8'd9;
    200: charMap = 8'd9;
    201: charMap = 8'd9;
    202: charMap = 8'd9;
    203: charMap = 8'd9;
    204: charMap = 8'd9;
    205: charMap = 8'd9;
    206: charMap = 8'd9;
    207: charMap = 8'd9;
    208: charMap = 8'd9;
    209: charMap = 8'd9;
    210: charMap = 8'd9;
    211: charMap = 8'd9;
    212: charMap = 8'd9;
    213: charMap = 8'd9;
    214: charMap = 8'd9;
    215: charMap = 8'd9;
    216: charMap = 8'd9;
    217: charMap = 8'd9;
    218: charMap = 8'd9;
    219: charMap = 8'd9;
    220: charMap = 8'd9;
    221: charMap = 8'd9;
    222: charMap = 8'd9;
    223: charMap = 8'd9;
    224: charMap = 8'd9;
    225: charMap = 8'd9;
    226: charMap = 8'd9;
    227: charMap = 8'd9;
    228: charMap = 8'd9;
    229: charMap = 8'd9;
    230: charMap = 8'd9;
    231: charMap = 8'd9;
    232: charMap = 8'd9;
    233: charMap = 8'd9;
    234: charMap = 8'd9;
    235: charMap = 8'd9;
    236: charMap = 8'd9;
    237: charMap = 8'd9;
    238: charMap = 8'd9;
    239: charMap = 8'd9;
    240: charMap = 8'd9;
    241: charMap = 8'd9;
    242: charMap = 8'd9;
    243: charMap = 8'd9;
    244: charMap = 8'd9;
    245: charMap = 8'd9;
    246: charMap = 8'd9;
    247: charMap = 8'd9;
    248: charMap = 8'd9;
    249: charMap = 8'd9;
    250: charMap = 8'd9;
    251: charMap = 8'd9;
    252: charMap = 8'd9;
    253: charMap = 8'd9;
    254: charMap = 8'd9;
    255: charMap = 8'd9;
    default: charMap = 8'bX;
  endcase
end
endfunction

function [10:0] stateMap;
  input [10:0] instate;
begin
  case( instate )
    0: stateMap = 11'd0;
    1: stateMap = 11'd1;
    2: stateMap = 11'd2;
    3: stateMap = 11'd3;
    4: stateMap = 11'd1;
    5: stateMap = 11'd4;
    6: stateMap = 11'd5;
    7: stateMap = 11'd6;
    8: stateMap = 11'd7;
    9: stateMap = 11'd8;
    10: stateMap = 11'd9;
    11: stateMap = 11'd10;
    12: stateMap = 11'd11;
    13: stateMap = 11'd12;
    14: stateMap = 11'd13;
    15: stateMap = 11'd14;
    16: stateMap = 11'd15;
    17: stateMap = 11'd16;
    18: stateMap = 11'd17;
    19: stateMap = 11'd18;
    20: stateMap = 11'd19;
    21: stateMap = 11'd20;
    22: stateMap = 11'd21;
    23: stateMap = 11'd22;
    24: stateMap = 11'd23;
    25: stateMap = 11'd24;
    26: stateMap = 11'd25;
    27: stateMap = 11'd26;
    28: stateMap = 11'd27;
    29: stateMap = 11'd28;
    30: stateMap = 11'd29;
    31: stateMap = 11'd30;
    32: stateMap = 11'd31;
    33: stateMap = 11'd32;
    34: stateMap = 11'd33;
    35: stateMap = 11'd34;
    36: stateMap = 11'd35;
    37: stateMap = 11'd36;
    38: stateMap = 11'd37;
    39: stateMap = 11'd38;
    40: stateMap = 11'd39;
    41: stateMap = 11'd40;
    42: stateMap = 11'd41;
    43: stateMap = 11'd42;
    44: stateMap = 11'd43;
    45: stateMap = 11'd44;
    46: stateMap = 11'd45;
    47: stateMap = 11'd46;
    48: stateMap = 11'd47;
    49: stateMap = 11'd48;
    50: stateMap = 11'd49;
    51: stateMap = 11'd50;
    52: stateMap = 11'd51;
    53: stateMap = 11'd2;
    54: stateMap = 11'd52;
    55: stateMap = 11'd2;
    56: stateMap = 11'd53;
    57: stateMap = 11'd54;
    58: stateMap = 11'd55;
    59: stateMap = 11'd56;
    60: stateMap = 11'd57;
    61: stateMap = 11'd58;
    62: stateMap = 11'd59;
    63: stateMap = 11'd60;
    64: stateMap = 11'd61;
    65: stateMap = 11'd62;
    66: stateMap = 11'd63;
    67: stateMap = 11'd64;
    68: stateMap = 11'd65;
    69: stateMap = 11'd66;
    70: stateMap = 11'd67;
    71: stateMap = 11'd68;
    72: stateMap = 11'd69;
    73: stateMap = 11'd70;
    74: stateMap = 11'd61;
    75: stateMap = 11'd71;
    76: stateMap = 11'd72;
    77: stateMap = 11'd73;
    78: stateMap = 11'd74;
    79: stateMap = 11'd75;
    80: stateMap = 11'd76;
    81: stateMap = 11'd77;
    82: stateMap = 11'd78;
    83: stateMap = 11'd79;
    84: stateMap = 11'd72;
    85: stateMap = 11'd80;
    86: stateMap = 11'd81;
    87: stateMap = 11'd82;
    88: stateMap = 11'd83;
    89: stateMap = 11'd84;
    90: stateMap = 11'd85;
    91: stateMap = 11'd86;
    92: stateMap = 11'd87;
    93: stateMap = 11'd88;
    94: stateMap = 11'd89;
    95: stateMap = 11'd90;
    96: stateMap = 11'd91;
    97: stateMap = 11'd92;
    98: stateMap = 11'd93;
    99: stateMap = 11'd83;
    100: stateMap = 11'd94;
    101: stateMap = 11'd95;
    102: stateMap = 11'd96;
    103: stateMap = 11'd97;
    104: stateMap = 11'd98;
    105: stateMap = 11'd99;
    106: stateMap = 11'd100;
    107: stateMap = 11'd101;
    108: stateMap = 11'd102;
    109: stateMap = 11'd103;
    110: stateMap = 11'd104;
    111: stateMap = 11'd105;
    112: stateMap = 11'd106;
    113: stateMap = 11'd107;
    114: stateMap = 11'd108;
    115: stateMap = 11'd109;
    116: stateMap = 11'd110;
    117: stateMap = 11'd111;
    118: stateMap = 11'd112;
    119: stateMap = 11'd113;
    120: stateMap = 11'd114;
    121: stateMap = 11'd115;
    122: stateMap = 11'd116;
    123: stateMap = 11'd117;
    124: stateMap = 11'd118;
    125: stateMap = 11'd119;
    126: stateMap = 11'd119;
    127: stateMap = 11'd120;
    128: stateMap = 11'd121;
    129: stateMap = 11'd122;
    130: stateMap = 11'd123;
    131: stateMap = 11'd124;
    132: stateMap = 11'd125;
    133: stateMap = 11'd126;
    134: stateMap = 11'd127;
    135: stateMap = 11'd128;
    136: stateMap = 11'd129;
    137: stateMap = 11'd130;
    138: stateMap = 11'd131;
    139: stateMap = 11'd132;
    140: stateMap = 11'd133;
    141: stateMap = 11'd134;
    142: stateMap = 11'd135;
    143: stateMap = 11'd136;
    144: stateMap = 11'd137;
    145: stateMap = 11'd123;
    146: stateMap = 11'd138;
    147: stateMap = 11'd139;
    148: stateMap = 11'd140;
    149: stateMap = 11'd141;
    150: stateMap = 11'd142;
    151: stateMap = 11'd143;
    152: stateMap = 11'd144;
    153: stateMap = 11'd145;
    154: stateMap = 11'd146;
    155: stateMap = 11'd147;
    156: stateMap = 11'd148;
    157: stateMap = 11'd149;
    158: stateMap = 11'd150;
    159: stateMap = 11'd151;
    160: stateMap = 11'd152;
    161: stateMap = 11'd153;
    162: stateMap = 11'd154;
    163: stateMap = 11'd155;
    164: stateMap = 11'd156;
    165: stateMap = 11'd157;
    166: stateMap = 11'd158;
    167: stateMap = 11'd159;
    168: stateMap = 11'd160;
    169: stateMap = 11'd161;
    170: stateMap = 11'd162;
    171: stateMap = 11'd163;
    172: stateMap = 11'd164;
    173: stateMap = 11'd165;
    174: stateMap = 11'd166;
    175: stateMap = 11'd167;
    176: stateMap = 11'd168;
    177: stateMap = 11'd169;
    178: stateMap = 11'd170;
    179: stateMap = 11'd171;
    180: stateMap = 11'd172;
    181: stateMap = 11'd173;
    182: stateMap = 11'd174;
    183: stateMap = 11'd175;
    184: stateMap = 11'd176;
    185: stateMap = 11'd177;
    186: stateMap = 11'd178;
    187: stateMap = 11'd179;
    188: stateMap = 11'd180;
    189: stateMap = 11'd181;
    190: stateMap = 11'd182;
    191: stateMap = 11'd183;
    192: stateMap = 11'd184;
    193: stateMap = 11'd185;
    194: stateMap = 11'd186;
    default: stateMap = 11'bX;
  endcase
end
endfunction

function acceptStates;
  input [10:0] instate;
begin
  case( instate )
    0: acceptStates = 1'b0;
    1: acceptStates = 1'b1;
    2: acceptStates = 1'b1;
    3: acceptStates = 1'b0;
    4: acceptStates = 1'b1;
    5: acceptStates = 1'b0;
    6: acceptStates = 1'b0;
    7: acceptStates = 1'b0;
    8: acceptStates = 1'b0;
    9: acceptStates = 1'b0;
    10: acceptStates = 1'b0;
    11: acceptStates = 1'b0;
    12: acceptStates = 1'b0;
    13: acceptStates = 1'b0;
    14: acceptStates = 1'b0;
    15: acceptStates = 1'b0;
    16: acceptStates = 1'b0;
    17: acceptStates = 1'b0;
    18: acceptStates = 1'b0;
    19: acceptStates = 1'b0;
    20: acceptStates = 1'b0;
    21: acceptStates = 1'b0;
    22: acceptStates = 1'b0;
    23: acceptStates = 1'b0;
    24: acceptStates = 1'b0;
    25: acceptStates = 1'b0;
    26: acceptStates = 1'b0;
    27: acceptStates = 1'b0;
    28: acceptStates = 1'b0;
    29: acceptStates = 1'b0;
    30: acceptStates = 1'b0;
    31: acceptStates = 1'b0;
    32: acceptStates = 1'b0;
    33: acceptStates = 1'b0;
    34: acceptStates = 1'b0;
    35: acceptStates = 1'b0;
    36: acceptStates = 1'b0;
    37: acceptStates = 1'b0;
    38: acceptStates = 1'b0;
    39: acceptStates = 1'b0;
    40: acceptStates = 1'b0;
    41: acceptStates = 1'b0;
    42: acceptStates = 1'b0;
    43: acceptStates = 1'b0;
    44: acceptStates = 1'b0;
    45: acceptStates = 1'b0;
    46: acceptStates = 1'b0;
    47: acceptStates = 1'b0;
    48: acceptStates = 1'b0;
    49: acceptStates = 1'b0;
    50: acceptStates = 1'b0;
    51: acceptStates = 1'b0;
    52: acceptStates = 1'b0;
    53: acceptStates = 1'b0;
    54: acceptStates = 1'b0;
    55: acceptStates = 1'b0;
    56: acceptStates = 1'b0;
    57: acceptStates = 1'b0;
    58: acceptStates = 1'b0;
    59: acceptStates = 1'b0;
    60: acceptStates = 1'b0;
    61: acceptStates = 1'b0;
    62: acceptStates = 1'b0;
    63: acceptStates = 1'b0;
    64: acceptStates = 1'b0;
    65: acceptStates = 1'b0;
    66: acceptStates = 1'b0;
    67: acceptStates = 1'b0;
    68: acceptStates = 1'b0;
    69: acceptStates = 1'b0;
    70: acceptStates = 1'b0;
    71: acceptStates = 1'b0;
    72: acceptStates = 1'b0;
    73: acceptStates = 1'b0;
    74: acceptStates = 1'b0;
    75: acceptStates = 1'b0;
    76: acceptStates = 1'b0;
    77: acceptStates = 1'b0;
    78: acceptStates = 1'b0;
    79: acceptStates = 1'b0;
    80: acceptStates = 1'b0;
    81: acceptStates = 1'b0;
    82: acceptStates = 1'b0;
    83: acceptStates = 1'b0;
    84: acceptStates = 1'b0;
    85: acceptStates = 1'b0;
    86: acceptStates = 1'b0;
    87: acceptStates = 1'b0;
    88: acceptStates = 1'b0;
    89: acceptStates = 1'b0;
    90: acceptStates = 1'b0;
    91: acceptStates = 1'b0;
    92: acceptStates = 1'b0;
    93: acceptStates = 1'b0;
    94: acceptStates = 1'b0;
    95: acceptStates = 1'b0;
    96: acceptStates = 1'b0;
    97: acceptStates = 1'b0;
    98: acceptStates = 1'b0;
    99: acceptStates = 1'b0;
    100: acceptStates = 1'b0;
    101: acceptStates = 1'b0;
    102: acceptStates = 1'b0;
    103: acceptStates = 1'b0;
    104: acceptStates = 1'b0;
    105: acceptStates = 1'b0;
    106: acceptStates = 1'b0;
    107: acceptStates = 1'b0;
    108: acceptStates = 1'b0;
    109: acceptStates = 1'b0;
    110: acceptStates = 1'b0;
    111: acceptStates = 1'b0;
    112: acceptStates = 1'b0;
    113: acceptStates = 1'b0;
    114: acceptStates = 1'b0;
    115: acceptStates = 1'b0;
    116: acceptStates = 1'b0;
    117: acceptStates = 1'b0;
    118: acceptStates = 1'b0;
    119: acceptStates = 1'b0;
    120: acceptStates = 1'b0;
    121: acceptStates = 1'b0;
    122: acceptStates = 1'b0;
    123: acceptStates = 1'b0;
    124: acceptStates = 1'b0;
    125: acceptStates = 1'b0;
    126: acceptStates = 1'b0;
    127: acceptStates = 1'b0;
    128: acceptStates = 1'b0;
    129: acceptStates = 1'b0;
    130: acceptStates = 1'b0;
    131: acceptStates = 1'b0;
    132: acceptStates = 1'b0;
    133: acceptStates = 1'b0;
    134: acceptStates = 1'b0;
    135: acceptStates = 1'b0;
    136: acceptStates = 1'b0;
    137: acceptStates = 1'b0;
    138: acceptStates = 1'b0;
    139: acceptStates = 1'b0;
    140: acceptStates = 1'b0;
    141: acceptStates = 1'b0;
    142: acceptStates = 1'b0;
    143: acceptStates = 1'b0;
    144: acceptStates = 1'b0;
    145: acceptStates = 1'b0;
    146: acceptStates = 1'b0;
    147: acceptStates = 1'b0;
    148: acceptStates = 1'b0;
    149: acceptStates = 1'b0;
    150: acceptStates = 1'b0;
    151: acceptStates = 1'b0;
    152: acceptStates = 1'b0;
    153: acceptStates = 1'b0;
    154: acceptStates = 1'b0;
    155: acceptStates = 1'b0;
    156: acceptStates = 1'b0;
    157: acceptStates = 1'b0;
    158: acceptStates = 1'b0;
    159: acceptStates = 1'b0;
    160: acceptStates = 1'b0;
    161: acceptStates = 1'b0;
    162: acceptStates = 1'b0;
    163: acceptStates = 1'b0;
    164: acceptStates = 1'b0;
    165: acceptStates = 1'b0;
    166: acceptStates = 1'b0;
    167: acceptStates = 1'b0;
    168: acceptStates = 1'b0;
    169: acceptStates = 1'b0;
    170: acceptStates = 1'b0;
    171: acceptStates = 1'b0;
    172: acceptStates = 1'b0;
    173: acceptStates = 1'b0;
    174: acceptStates = 1'b0;
    175: acceptStates = 1'b0;
    176: acceptStates = 1'b0;
    177: acceptStates = 1'b0;
    178: acceptStates = 1'b0;
    179: acceptStates = 1'b0;
    180: acceptStates = 1'b0;
    181: acceptStates = 1'b0;
    182: acceptStates = 1'b0;
    183: acceptStates = 1'b0;
    184: acceptStates = 1'b0;
    185: acceptStates = 1'b0;
    186: acceptStates = 1'b0;
    187: acceptStates = 1'b0;
    188: acceptStates = 1'b0;
    189: acceptStates = 1'b0;
    190: acceptStates = 1'b0;
    191: acceptStates = 1'b0;
    192: acceptStates = 1'b0;
    193: acceptStates = 1'b0;
    194: acceptStates = 1'b0;
    default: acceptStates = 1'bX;
  endcase
end
endfunction

function [10:0] stateTransition;
  input [10:0] mapped_state;
  input [7:0]  mapped_char;
begin
  case( mapped_state )
    0: case ( mapped_char ) 
      0: stateTransition = 11'd1;
      1: stateTransition = 11'd3;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    1: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    2: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    3: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd5;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    4: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd6;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    5: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd7;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    6: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd8;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    7: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd9;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    8: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd10;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    9: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd11;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    10: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd12;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    11: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd13;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    12: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd14;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    13: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd15;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    14: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd16;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    15: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd17;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    16: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd18;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    17: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    18: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    19: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd20;
      22: stateTransition = 11'd21;
      23: stateTransition = 11'd22;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    20: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd21;
      22: stateTransition = 11'd21;
      23: stateTransition = 11'd23;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    21: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd2;
      25: stateTransition = 11'd2;
      26: stateTransition = 11'd39;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd24;
      default: stateTransition = 11'bX;
    endcase
    22: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd4;
      25: stateTransition = 11'd4;
      26: stateTransition = 11'd25;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd26;
      default: stateTransition = 11'bX;
    endcase
    23: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd2;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    24: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd27;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    25: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd4;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    26: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd28;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    27: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd29;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    28: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd31;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd0;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    29: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd2;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    30: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd0;
      2: stateTransition = 11'd0;
      3: stateTransition = 11'd0;
      4: stateTransition = 11'd0;
      5: stateTransition = 11'd0;
      6: stateTransition = 11'd0;
      7: stateTransition = 11'd0;
      8: stateTransition = 11'd0;
      9: stateTransition = 11'd0;
      10: stateTransition = 11'd0;
      11: stateTransition = 11'd0;
      12: stateTransition = 11'd0;
      13: stateTransition = 11'd0;
      14: stateTransition = 11'd0;
      15: stateTransition = 11'd0;
      16: stateTransition = 11'd0;
      17: stateTransition = 11'd0;
      18: stateTransition = 11'd0;
      19: stateTransition = 11'd0;
      20: stateTransition = 11'd0;
      21: stateTransition = 11'd0;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd0;
      24: stateTransition = 11'd0;
      25: stateTransition = 11'd0;
      26: stateTransition = 11'd0;
      27: stateTransition = 11'd0;
      28: stateTransition = 11'd4;
      29: stateTransition = 11'd0;
      default: stateTransition = 11'bX;
    endcase
    31: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd20;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    32: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd30;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    33: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd32;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    34: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd50;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd33;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    35: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd34;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    36: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd35;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    37: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd36;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    38: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd37;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    39: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd38;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    40: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd40;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    41: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd41;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    42: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd42;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd110;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd147;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    43: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd43;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    44: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd44;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    45: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd45;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    46: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd46;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    47: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd47;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    48: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd48;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd194;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    49: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd48;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    50: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd49;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    51: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd50;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    52: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd51;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd161;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    53: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd54;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    54: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    55: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd132;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd56;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    56: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd55;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    57: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd56;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    58: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd57;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd131;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    59: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd58;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    60: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd57;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    61: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd62;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    62: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd57;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    63: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd57;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd131;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    64: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd72;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    65: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd57;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    66: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd111;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd127;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd129;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    67: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd98;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd59;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    68: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd60;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    69: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd74;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    70: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd61;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    71: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd63;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    72: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd71;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    73: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd65;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    74: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd64;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    75: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd66;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    76: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd67;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    77: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd68;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    78: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd69;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    79: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd70;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    80: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd176;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd73;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    81: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd76;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    82: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd75;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    83: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd86;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    84: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd77;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    85: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd78;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    86: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd79;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    87: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd74;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    88: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd80;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    89: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd81;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    90: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd82;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd166;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    91: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd83;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd129;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    92: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd84;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    93: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd85;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    94: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd87;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    95: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd88;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    96: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd89;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    97: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd90;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    98: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd91;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    99: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd92;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    100: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd93;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    101: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd94;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    102: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd95;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    103: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd96;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    104: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd99;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    105: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    106: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd98;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    107: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd101;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd147;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    108: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd189;
      5: stateTransition = 11'd109;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    109: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd136;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd110;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd147;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    110: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd100;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    111: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd103;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    112: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd102;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    113: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd105;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    114: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd104;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    115: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd106;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd131;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    116: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd107;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    117: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd108;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    118: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd109;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    119: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd110;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd147;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    120: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd112;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    121: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd113;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    122: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd114;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    123: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd128;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    124: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd116;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    125: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd115;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    126: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd118;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    127: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd117;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    128: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd165;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd131;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    129: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd126;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    130: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd120;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    131: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd119;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    132: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd121;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    133: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd122;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    134: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd123;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    135: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd124;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    136: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd125;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    137: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd127;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd129;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    138: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd131;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    139: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd130;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    140: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd133;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    141: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd134;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    142: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd135;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    143: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd138;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    144: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd137;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    145: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd191;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd139;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    146: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd140;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    147: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd141;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    148: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd144;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    149: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd145;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    150: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd181;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd131;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    151: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd158;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    152: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd146;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    153: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd149;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    154: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd148;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    155: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd151;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    156: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd150;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    157: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd152;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    158: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd153;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    159: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd154;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    160: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd159;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    161: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd155;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    162: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd164;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    163: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd163;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    164: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd166;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    165: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd167;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    166: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd168;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    167: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd169;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    168: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd172;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    169: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd171;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    170: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd173;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    171: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd186;
      4: stateTransition = 11'd176;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    172: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd174;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    173: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd175;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    174: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd176;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    175: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd177;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    176: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd178;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    177: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd179;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    178: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd180;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    179: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd182;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    180: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd183;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    181: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd184;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    182: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd19;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd185;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    183: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd19;
      2: stateTransition = 11'd190;
      3: stateTransition = 11'd19;
      4: stateTransition = 11'd19;
      5: stateTransition = 11'd156;
      6: stateTransition = 11'd19;
      7: stateTransition = 11'd160;
      8: stateTransition = 11'd170;
      9: stateTransition = 11'd19;
      10: stateTransition = 11'd187;
      11: stateTransition = 11'd19;
      12: stateTransition = 11'd19;
      13: stateTransition = 11'd19;
      14: stateTransition = 11'd19;
      15: stateTransition = 11'd19;
      16: stateTransition = 11'd19;
      17: stateTransition = 11'd142;
      18: stateTransition = 11'd162;
      19: stateTransition = 11'd19;
      20: stateTransition = 11'd19;
      21: stateTransition = 11'd19;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd19;
      24: stateTransition = 11'd19;
      25: stateTransition = 11'd19;
      26: stateTransition = 11'd19;
      27: stateTransition = 11'd19;
      28: stateTransition = 11'd19;
      29: stateTransition = 11'd19;
      default: stateTransition = 11'bX;
    endcase
    184: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd188;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    185: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd53;
      3: stateTransition = 11'd192;
      4: stateTransition = 11'd71;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    186: case ( mapped_char ) 
      0: stateTransition = 11'd0;
      1: stateTransition = 11'd52;
      2: stateTransition = 11'd193;
      3: stateTransition = 11'd53;
      4: stateTransition = 11'd53;
      5: stateTransition = 11'd143;
      6: stateTransition = 11'd53;
      7: stateTransition = 11'd53;
      8: stateTransition = 11'd53;
      9: stateTransition = 11'd53;
      10: stateTransition = 11'd97;
      11: stateTransition = 11'd53;
      12: stateTransition = 11'd53;
      13: stateTransition = 11'd53;
      14: stateTransition = 11'd53;
      15: stateTransition = 11'd53;
      16: stateTransition = 11'd53;
      17: stateTransition = 11'd157;
      18: stateTransition = 11'd53;
      19: stateTransition = 11'd53;
      20: stateTransition = 11'd53;
      21: stateTransition = 11'd53;
      22: stateTransition = 11'd0;
      23: stateTransition = 11'd53;
      24: stateTransition = 11'd53;
      25: stateTransition = 11'd53;
      26: stateTransition = 11'd53;
      27: stateTransition = 11'd53;
      28: stateTransition = 11'd53;
      29: stateTransition = 11'd53;
      default: stateTransition = 11'bX;
    endcase
    default: stateTransition = 11'bX;
  endcase
end
endfunction

`else

function [7:0] charMap;
input [7:0] inchar;
begin
    charMap = inchar;
end
endfunction

function [10:0] stateMap;
input [10:0] instate;
begin
    stateMap = instate;
end
endfunction

function acceptStates;
    input [10:0] instate;
begin
    acceptStates = 1'b0;
end
endfunction

function [10:0] stateTransition;
    input [10:0] instate;
    input [7:0]  inchar;
begin
    stateTransition = instate;
end
endfunction

`endif

    // Invoke the DFA functions.
    wire [7:0]  mapped_char;
    wire [10:0] mapped_state, next_state;
    wire next_accept;
    assign mapped_char = charMap(char_in);
    assign mapped_state = stateMap(cur_state);
    assign next_state = stateTransition(mapped_state, mapped_char);
    assign next_accept = acceptStates(next_state);
    // Update our outputs.
    assign accept_out = state_in_vld ? 1'b0 : char_in_vld ? next_accept : 1'b0;
    assign state_out = cur_state;
    // Update our local state.
    always @(posedge clk)
    begin
       if (!rst_n)
        begin
            cur_state <= 0;
        end
        else
        begin
            if (state_in_vld)
            begin
                cur_state <= state_in;
            end
            else if (char_in_vld)
            begin
                cur_state <= next_state;
            end
        end
    end
endmodule
