wire [15:0] count_ALL_0 ;
wire [15:0] count_ALL_1 ;
wire [15:0] count_ALL_2 ;
wire [15:0] count_ALL_3 ;
wire [15:0] count_ALL_4 ;
wire [15:0] count_finger_0 ;
wire [15:0] count_ftp_0 ;
wire [15:0] count_http_0 ;
wire [15:0] count_imap_0 ;
wire [15:0] count_netbios_0 ;
wire [15:0] count_nntp_0 ;
wire [15:0] count_pop3_0 ;
wire [15:0] count_rlogin_0 ;
wire [15:0] count_smtp_0 ;
wire [15:0] count_telnet_0 ;
wire [15:0] count_CATEGORY_finger ;
wire [15:0] count_CATEGORY_ftp ;
wire [15:0] count_CATEGORY_http ;
wire [15:0] count_CATEGORY_imap ;
wire [15:0] count_CATEGORY_netbios ;
wire [15:0] count_CATEGORY_nntp ;
wire [15:0] count_CATEGORY_pop3 ;
wire [15:0] count_CATEGORY_rlogin ;
wire [15:0] count_CATEGORY_smtp ;
wire [15:0] count_CATEGORY_telnet ;

`ifdef REGEX_OPTIONAL
wire [15:0] count_ALL_5 ;
wire [15:0] count_ALL_6 ;
wire [15:0] count_ALL_7 ;
wire [15:0] count_ALL_8 ;
wire [15:0] count_ALL_9 ;
wire [15:0] count_ALL_10 ;
wire [15:0] count_ALL_11 ;
wire [15:0] count_ALL_12 ;
wire [15:0] count_ALL_13 ;
wire [15:0] count_ALL_14 ;



wire [15:0] count_finger_1 ;
wire [15:0] count_finger_2 ;
wire [15:0] count_finger_3 ;
wire [15:0] count_finger_4 ;
wire [15:0] count_finger_5 ;

wire [15:0] count_ftp_1 ;
wire [15:0] count_ftp_2 ;
wire [15:0] count_ftp_3 ;
wire [15:0] count_ftp_4 ;
wire [15:0] count_ftp_5 ;
wire [15:0] count_ftp_6 ;
wire [15:0] count_ftp_7 ;
wire [15:0] count_ftp_8 ;
wire [15:0] count_ftp_9 ;



wire [15:0] count_http_1 ;
wire [15:0] count_http_2 ;
wire [15:0] count_http_3 ;
wire [15:0] count_http_4 ;
wire [15:0] count_http_5 ;
wire [15:0] count_http_6 ;
wire [15:0] count_http_7 ;
wire [15:0] count_http_8 ;
wire [15:0] count_http_9 ;

wire [15:0] count_imap_1 ;
wire [15:0] count_imap_2 ;
wire [15:0] count_imap_3 ;
wire [15:0] count_imap_4 ;
wire [15:0] count_imap_5 ;
wire [15:0] count_imap_6 ;
wire [15:0] count_imap_7 ;
wire [15:0] count_imap_8 ;
wire [15:0] count_imap_9 ;

wire [15:0] count_netbios_1 ;
wire [15:0] count_netbios_2 ;
wire [15:0] count_netbios_3 ;
wire [15:0] count_netbios_4 ;
wire [15:0] count_netbios_5 ;
wire [15:0] count_netbios_6 ;
wire [15:0] count_netbios_7 ;
wire [15:0] count_netbios_8 ;
wire [15:0] count_netbios_9 ;

wire [15:0] count_nntp_1 ;
wire [15:0] count_nntp_2 ;
wire [15:0] count_nntp_3 ;
wire [15:0] count_nntp_4 ;
wire [15:0] count_nntp_5 ;
wire [15:0] count_nntp_6 ;
wire [15:0] count_nntp_7 ;
wire [15:0] count_nntp_8 ;
wire [15:0] count_nntp_9 ;

wire [15:0] count_pop3_1 ;
wire [15:0] count_pop3_2 ;
wire [15:0] count_pop3_3 ;
wire [15:0] count_pop3_4 ;
wire [15:0] count_pop3_5 ;
wire [15:0] count_pop3_6 ;
wire [15:0] count_pop3_7 ;
wire [15:0] count_pop3_8 ;
wire [15:0] count_pop3_9 ;


wire [15:0] count_rlogin_1 ;
wire [15:0] count_rlogin_2 ;
wire [15:0] count_rlogin_3 ;
wire [15:0] count_rlogin_4 ;
wire [15:0] count_rlogin_5 ;


wire [15:0] count_smtp_1 ;
wire [15:0] count_smtp_2 ;
wire [15:0] count_smtp_3 ;
wire [15:0] count_smtp_4 ;
wire [15:0] count_smtp_5 ;
wire [15:0] count_smtp_6 ;
wire [15:0] count_smtp_7 ;
wire [15:0] count_smtp_8 ;
wire [15:0] count_smtp_9 ;


wire [15:0] count_telnet_1 ;
wire [15:0] count_telnet_2 ;
wire [15:0] count_telnet_3 ;
wire [15:0] count_telnet_4 ;
wire [15:0] count_telnet_5 ;
wire [15:0] count_telnet_6 ;
wire [15:0] count_telnet_7 ;
wire [15:0] count_telnet_8 ;
wire [15:0] count_telnet_9 ;

wire [15:0] count_CATEGORY_aim ;
wire [15:0] count_CATEGORY_bittorrent ;
wire [15:0] count_CATEGORY_cvs ;
wire [15:0] count_CATEGORY_dhcp ;
wire [15:0] count_CATEGORY_directconnect ;
wire [15:0] count_CATEGORY_dns ;
wire [15:0] count_CATEGORY_fasttrack ;
wire [15:0] count_CATEGORY_tor ;
wire [15:0] count_CATEGORY_vnc ;
wire [15:0] count_CATEGORY_worldofwarcraft ;
wire [15:0] count_CATEGORY_x11 ;
wire [15:0] count_CATEGORY_yahoo ;
wire [15:0] count_CATEGORY_freenet ;
wire [15:0] count_CATEGORY_gnutella ;
wire [15:0] count_CATEGORY_gopher ;
wire [15:0] count_CATEGORY_irc ;
wire [15:0] count_CATEGORY_jabber ;
wire [15:0] count_CATEGORY_msn ;
wire [15:0] count_CATEGORY_napster ;
wire [15:0] count_CATEGORY_sip ;
wire [15:0] count_CATEGORY_snmp ;
wire [15:0] count_CATEGORY_socks ;
wire [15:0] count_CATEGORY_ssh ;
wire [15:0] count_CATEGORY_ssl ;
wire [15:0] count_CATEGORY_subversion ;
`endif //  `ifdef REGEX_OPTIONAL
