module tb;

   tag_parser dut_i (/*AUTOINST*/);
   
   
endmodule // tb
